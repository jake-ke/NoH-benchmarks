`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO = "Knn_Knn,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvh1582-vsva3697-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=3956,HLS_SYN_LUT=7208,HLS_VERSION=2023_2_2}" *)


module Knn
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_L4_out_dist_ARADDR,
  m_axi_L4_out_dist_ARBURST,
  m_axi_L4_out_dist_ARCACHE,
  m_axi_L4_out_dist_ARID,
  m_axi_L4_out_dist_ARLEN,
  m_axi_L4_out_dist_ARLOCK,
  m_axi_L4_out_dist_ARPROT,
  m_axi_L4_out_dist_ARQOS,
  m_axi_L4_out_dist_ARREADY,
  m_axi_L4_out_dist_ARSIZE,
  m_axi_L4_out_dist_ARVALID,
  m_axi_L4_out_dist_AWADDR,
  m_axi_L4_out_dist_AWBURST,
  m_axi_L4_out_dist_AWCACHE,
  m_axi_L4_out_dist_AWID,
  m_axi_L4_out_dist_AWLEN,
  m_axi_L4_out_dist_AWLOCK,
  m_axi_L4_out_dist_AWPROT,
  m_axi_L4_out_dist_AWQOS,
  m_axi_L4_out_dist_AWREADY,
  m_axi_L4_out_dist_AWSIZE,
  m_axi_L4_out_dist_AWVALID,
  m_axi_L4_out_dist_BID,
  m_axi_L4_out_dist_BREADY,
  m_axi_L4_out_dist_BRESP,
  m_axi_L4_out_dist_BVALID,
  m_axi_L4_out_dist_RDATA,
  m_axi_L4_out_dist_RID,
  m_axi_L4_out_dist_RLAST,
  m_axi_L4_out_dist_RREADY,
  m_axi_L4_out_dist_RRESP,
  m_axi_L4_out_dist_RVALID,
  m_axi_L4_out_dist_WDATA,
  m_axi_L4_out_dist_WLAST,
  m_axi_L4_out_dist_WREADY,
  m_axi_L4_out_dist_WSTRB,
  m_axi_L4_out_dist_WVALID,
  m_axi_L4_out_id_ARADDR,
  m_axi_L4_out_id_ARBURST,
  m_axi_L4_out_id_ARCACHE,
  m_axi_L4_out_id_ARID,
  m_axi_L4_out_id_ARLEN,
  m_axi_L4_out_id_ARLOCK,
  m_axi_L4_out_id_ARPROT,
  m_axi_L4_out_id_ARQOS,
  m_axi_L4_out_id_ARREADY,
  m_axi_L4_out_id_ARSIZE,
  m_axi_L4_out_id_ARVALID,
  m_axi_L4_out_id_AWADDR,
  m_axi_L4_out_id_AWBURST,
  m_axi_L4_out_id_AWCACHE,
  m_axi_L4_out_id_AWID,
  m_axi_L4_out_id_AWLEN,
  m_axi_L4_out_id_AWLOCK,
  m_axi_L4_out_id_AWPROT,
  m_axi_L4_out_id_AWQOS,
  m_axi_L4_out_id_AWREADY,
  m_axi_L4_out_id_AWSIZE,
  m_axi_L4_out_id_AWVALID,
  m_axi_L4_out_id_BID,
  m_axi_L4_out_id_BREADY,
  m_axi_L4_out_id_BRESP,
  m_axi_L4_out_id_BVALID,
  m_axi_L4_out_id_RDATA,
  m_axi_L4_out_id_RID,
  m_axi_L4_out_id_RLAST,
  m_axi_L4_out_id_RREADY,
  m_axi_L4_out_id_RRESP,
  m_axi_L4_out_id_RVALID,
  m_axi_L4_out_id_WDATA,
  m_axi_L4_out_id_WLAST,
  m_axi_L4_out_id_WREADY,
  m_axi_L4_out_id_WSTRB,
  m_axi_L4_out_id_WVALID,
  m_axi_in_0_ARADDR,
  m_axi_in_0_ARBURST,
  m_axi_in_0_ARCACHE,
  m_axi_in_0_ARID,
  m_axi_in_0_ARLEN,
  m_axi_in_0_ARLOCK,
  m_axi_in_0_ARPROT,
  m_axi_in_0_ARQOS,
  m_axi_in_0_ARREADY,
  m_axi_in_0_ARSIZE,
  m_axi_in_0_ARVALID,
  m_axi_in_0_AWADDR,
  m_axi_in_0_AWBURST,
  m_axi_in_0_AWCACHE,
  m_axi_in_0_AWID,
  m_axi_in_0_AWLEN,
  m_axi_in_0_AWLOCK,
  m_axi_in_0_AWPROT,
  m_axi_in_0_AWQOS,
  m_axi_in_0_AWREADY,
  m_axi_in_0_AWSIZE,
  m_axi_in_0_AWVALID,
  m_axi_in_0_BID,
  m_axi_in_0_BREADY,
  m_axi_in_0_BRESP,
  m_axi_in_0_BVALID,
  m_axi_in_0_RDATA,
  m_axi_in_0_RID,
  m_axi_in_0_RLAST,
  m_axi_in_0_RREADY,
  m_axi_in_0_RRESP,
  m_axi_in_0_RVALID,
  m_axi_in_0_WDATA,
  m_axi_in_0_WLAST,
  m_axi_in_0_WREADY,
  m_axi_in_0_WSTRB,
  m_axi_in_0_WVALID,
  m_axi_in_1_ARADDR,
  m_axi_in_1_ARBURST,
  m_axi_in_1_ARCACHE,
  m_axi_in_1_ARID,
  m_axi_in_1_ARLEN,
  m_axi_in_1_ARLOCK,
  m_axi_in_1_ARPROT,
  m_axi_in_1_ARQOS,
  m_axi_in_1_ARREADY,
  m_axi_in_1_ARSIZE,
  m_axi_in_1_ARVALID,
  m_axi_in_1_AWADDR,
  m_axi_in_1_AWBURST,
  m_axi_in_1_AWCACHE,
  m_axi_in_1_AWID,
  m_axi_in_1_AWLEN,
  m_axi_in_1_AWLOCK,
  m_axi_in_1_AWPROT,
  m_axi_in_1_AWQOS,
  m_axi_in_1_AWREADY,
  m_axi_in_1_AWSIZE,
  m_axi_in_1_AWVALID,
  m_axi_in_1_BID,
  m_axi_in_1_BREADY,
  m_axi_in_1_BRESP,
  m_axi_in_1_BVALID,
  m_axi_in_1_RDATA,
  m_axi_in_1_RID,
  m_axi_in_1_RLAST,
  m_axi_in_1_RREADY,
  m_axi_in_1_RRESP,
  m_axi_in_1_RVALID,
  m_axi_in_1_WDATA,
  m_axi_in_1_WLAST,
  m_axi_in_1_WREADY,
  m_axi_in_1_WSTRB,
  m_axi_in_1_WVALID,
  m_axi_in_10_ARADDR,
  m_axi_in_10_ARBURST,
  m_axi_in_10_ARCACHE,
  m_axi_in_10_ARID,
  m_axi_in_10_ARLEN,
  m_axi_in_10_ARLOCK,
  m_axi_in_10_ARPROT,
  m_axi_in_10_ARQOS,
  m_axi_in_10_ARREADY,
  m_axi_in_10_ARSIZE,
  m_axi_in_10_ARVALID,
  m_axi_in_10_AWADDR,
  m_axi_in_10_AWBURST,
  m_axi_in_10_AWCACHE,
  m_axi_in_10_AWID,
  m_axi_in_10_AWLEN,
  m_axi_in_10_AWLOCK,
  m_axi_in_10_AWPROT,
  m_axi_in_10_AWQOS,
  m_axi_in_10_AWREADY,
  m_axi_in_10_AWSIZE,
  m_axi_in_10_AWVALID,
  m_axi_in_10_BID,
  m_axi_in_10_BREADY,
  m_axi_in_10_BRESP,
  m_axi_in_10_BVALID,
  m_axi_in_10_RDATA,
  m_axi_in_10_RID,
  m_axi_in_10_RLAST,
  m_axi_in_10_RREADY,
  m_axi_in_10_RRESP,
  m_axi_in_10_RVALID,
  m_axi_in_10_WDATA,
  m_axi_in_10_WLAST,
  m_axi_in_10_WREADY,
  m_axi_in_10_WSTRB,
  m_axi_in_10_WVALID,
  m_axi_in_11_ARADDR,
  m_axi_in_11_ARBURST,
  m_axi_in_11_ARCACHE,
  m_axi_in_11_ARID,
  m_axi_in_11_ARLEN,
  m_axi_in_11_ARLOCK,
  m_axi_in_11_ARPROT,
  m_axi_in_11_ARQOS,
  m_axi_in_11_ARREADY,
  m_axi_in_11_ARSIZE,
  m_axi_in_11_ARVALID,
  m_axi_in_11_AWADDR,
  m_axi_in_11_AWBURST,
  m_axi_in_11_AWCACHE,
  m_axi_in_11_AWID,
  m_axi_in_11_AWLEN,
  m_axi_in_11_AWLOCK,
  m_axi_in_11_AWPROT,
  m_axi_in_11_AWQOS,
  m_axi_in_11_AWREADY,
  m_axi_in_11_AWSIZE,
  m_axi_in_11_AWVALID,
  m_axi_in_11_BID,
  m_axi_in_11_BREADY,
  m_axi_in_11_BRESP,
  m_axi_in_11_BVALID,
  m_axi_in_11_RDATA,
  m_axi_in_11_RID,
  m_axi_in_11_RLAST,
  m_axi_in_11_RREADY,
  m_axi_in_11_RRESP,
  m_axi_in_11_RVALID,
  m_axi_in_11_WDATA,
  m_axi_in_11_WLAST,
  m_axi_in_11_WREADY,
  m_axi_in_11_WSTRB,
  m_axi_in_11_WVALID,
  m_axi_in_12_ARADDR,
  m_axi_in_12_ARBURST,
  m_axi_in_12_ARCACHE,
  m_axi_in_12_ARID,
  m_axi_in_12_ARLEN,
  m_axi_in_12_ARLOCK,
  m_axi_in_12_ARPROT,
  m_axi_in_12_ARQOS,
  m_axi_in_12_ARREADY,
  m_axi_in_12_ARSIZE,
  m_axi_in_12_ARVALID,
  m_axi_in_12_AWADDR,
  m_axi_in_12_AWBURST,
  m_axi_in_12_AWCACHE,
  m_axi_in_12_AWID,
  m_axi_in_12_AWLEN,
  m_axi_in_12_AWLOCK,
  m_axi_in_12_AWPROT,
  m_axi_in_12_AWQOS,
  m_axi_in_12_AWREADY,
  m_axi_in_12_AWSIZE,
  m_axi_in_12_AWVALID,
  m_axi_in_12_BID,
  m_axi_in_12_BREADY,
  m_axi_in_12_BRESP,
  m_axi_in_12_BVALID,
  m_axi_in_12_RDATA,
  m_axi_in_12_RID,
  m_axi_in_12_RLAST,
  m_axi_in_12_RREADY,
  m_axi_in_12_RRESP,
  m_axi_in_12_RVALID,
  m_axi_in_12_WDATA,
  m_axi_in_12_WLAST,
  m_axi_in_12_WREADY,
  m_axi_in_12_WSTRB,
  m_axi_in_12_WVALID,
  m_axi_in_13_ARADDR,
  m_axi_in_13_ARBURST,
  m_axi_in_13_ARCACHE,
  m_axi_in_13_ARID,
  m_axi_in_13_ARLEN,
  m_axi_in_13_ARLOCK,
  m_axi_in_13_ARPROT,
  m_axi_in_13_ARQOS,
  m_axi_in_13_ARREADY,
  m_axi_in_13_ARSIZE,
  m_axi_in_13_ARVALID,
  m_axi_in_13_AWADDR,
  m_axi_in_13_AWBURST,
  m_axi_in_13_AWCACHE,
  m_axi_in_13_AWID,
  m_axi_in_13_AWLEN,
  m_axi_in_13_AWLOCK,
  m_axi_in_13_AWPROT,
  m_axi_in_13_AWQOS,
  m_axi_in_13_AWREADY,
  m_axi_in_13_AWSIZE,
  m_axi_in_13_AWVALID,
  m_axi_in_13_BID,
  m_axi_in_13_BREADY,
  m_axi_in_13_BRESP,
  m_axi_in_13_BVALID,
  m_axi_in_13_RDATA,
  m_axi_in_13_RID,
  m_axi_in_13_RLAST,
  m_axi_in_13_RREADY,
  m_axi_in_13_RRESP,
  m_axi_in_13_RVALID,
  m_axi_in_13_WDATA,
  m_axi_in_13_WLAST,
  m_axi_in_13_WREADY,
  m_axi_in_13_WSTRB,
  m_axi_in_13_WVALID,
  m_axi_in_14_ARADDR,
  m_axi_in_14_ARBURST,
  m_axi_in_14_ARCACHE,
  m_axi_in_14_ARID,
  m_axi_in_14_ARLEN,
  m_axi_in_14_ARLOCK,
  m_axi_in_14_ARPROT,
  m_axi_in_14_ARQOS,
  m_axi_in_14_ARREADY,
  m_axi_in_14_ARSIZE,
  m_axi_in_14_ARVALID,
  m_axi_in_14_AWADDR,
  m_axi_in_14_AWBURST,
  m_axi_in_14_AWCACHE,
  m_axi_in_14_AWID,
  m_axi_in_14_AWLEN,
  m_axi_in_14_AWLOCK,
  m_axi_in_14_AWPROT,
  m_axi_in_14_AWQOS,
  m_axi_in_14_AWREADY,
  m_axi_in_14_AWSIZE,
  m_axi_in_14_AWVALID,
  m_axi_in_14_BID,
  m_axi_in_14_BREADY,
  m_axi_in_14_BRESP,
  m_axi_in_14_BVALID,
  m_axi_in_14_RDATA,
  m_axi_in_14_RID,
  m_axi_in_14_RLAST,
  m_axi_in_14_RREADY,
  m_axi_in_14_RRESP,
  m_axi_in_14_RVALID,
  m_axi_in_14_WDATA,
  m_axi_in_14_WLAST,
  m_axi_in_14_WREADY,
  m_axi_in_14_WSTRB,
  m_axi_in_14_WVALID,
  m_axi_in_15_ARADDR,
  m_axi_in_15_ARBURST,
  m_axi_in_15_ARCACHE,
  m_axi_in_15_ARID,
  m_axi_in_15_ARLEN,
  m_axi_in_15_ARLOCK,
  m_axi_in_15_ARPROT,
  m_axi_in_15_ARQOS,
  m_axi_in_15_ARREADY,
  m_axi_in_15_ARSIZE,
  m_axi_in_15_ARVALID,
  m_axi_in_15_AWADDR,
  m_axi_in_15_AWBURST,
  m_axi_in_15_AWCACHE,
  m_axi_in_15_AWID,
  m_axi_in_15_AWLEN,
  m_axi_in_15_AWLOCK,
  m_axi_in_15_AWPROT,
  m_axi_in_15_AWQOS,
  m_axi_in_15_AWREADY,
  m_axi_in_15_AWSIZE,
  m_axi_in_15_AWVALID,
  m_axi_in_15_BID,
  m_axi_in_15_BREADY,
  m_axi_in_15_BRESP,
  m_axi_in_15_BVALID,
  m_axi_in_15_RDATA,
  m_axi_in_15_RID,
  m_axi_in_15_RLAST,
  m_axi_in_15_RREADY,
  m_axi_in_15_RRESP,
  m_axi_in_15_RVALID,
  m_axi_in_15_WDATA,
  m_axi_in_15_WLAST,
  m_axi_in_15_WREADY,
  m_axi_in_15_WSTRB,
  m_axi_in_15_WVALID,
  m_axi_in_16_ARADDR,
  m_axi_in_16_ARBURST,
  m_axi_in_16_ARCACHE,
  m_axi_in_16_ARID,
  m_axi_in_16_ARLEN,
  m_axi_in_16_ARLOCK,
  m_axi_in_16_ARPROT,
  m_axi_in_16_ARQOS,
  m_axi_in_16_ARREADY,
  m_axi_in_16_ARSIZE,
  m_axi_in_16_ARVALID,
  m_axi_in_16_AWADDR,
  m_axi_in_16_AWBURST,
  m_axi_in_16_AWCACHE,
  m_axi_in_16_AWID,
  m_axi_in_16_AWLEN,
  m_axi_in_16_AWLOCK,
  m_axi_in_16_AWPROT,
  m_axi_in_16_AWQOS,
  m_axi_in_16_AWREADY,
  m_axi_in_16_AWSIZE,
  m_axi_in_16_AWVALID,
  m_axi_in_16_BID,
  m_axi_in_16_BREADY,
  m_axi_in_16_BRESP,
  m_axi_in_16_BVALID,
  m_axi_in_16_RDATA,
  m_axi_in_16_RID,
  m_axi_in_16_RLAST,
  m_axi_in_16_RREADY,
  m_axi_in_16_RRESP,
  m_axi_in_16_RVALID,
  m_axi_in_16_WDATA,
  m_axi_in_16_WLAST,
  m_axi_in_16_WREADY,
  m_axi_in_16_WSTRB,
  m_axi_in_16_WVALID,
  m_axi_in_17_ARADDR,
  m_axi_in_17_ARBURST,
  m_axi_in_17_ARCACHE,
  m_axi_in_17_ARID,
  m_axi_in_17_ARLEN,
  m_axi_in_17_ARLOCK,
  m_axi_in_17_ARPROT,
  m_axi_in_17_ARQOS,
  m_axi_in_17_ARREADY,
  m_axi_in_17_ARSIZE,
  m_axi_in_17_ARVALID,
  m_axi_in_17_AWADDR,
  m_axi_in_17_AWBURST,
  m_axi_in_17_AWCACHE,
  m_axi_in_17_AWID,
  m_axi_in_17_AWLEN,
  m_axi_in_17_AWLOCK,
  m_axi_in_17_AWPROT,
  m_axi_in_17_AWQOS,
  m_axi_in_17_AWREADY,
  m_axi_in_17_AWSIZE,
  m_axi_in_17_AWVALID,
  m_axi_in_17_BID,
  m_axi_in_17_BREADY,
  m_axi_in_17_BRESP,
  m_axi_in_17_BVALID,
  m_axi_in_17_RDATA,
  m_axi_in_17_RID,
  m_axi_in_17_RLAST,
  m_axi_in_17_RREADY,
  m_axi_in_17_RRESP,
  m_axi_in_17_RVALID,
  m_axi_in_17_WDATA,
  m_axi_in_17_WLAST,
  m_axi_in_17_WREADY,
  m_axi_in_17_WSTRB,
  m_axi_in_17_WVALID,
  m_axi_in_18_ARADDR,
  m_axi_in_18_ARBURST,
  m_axi_in_18_ARCACHE,
  m_axi_in_18_ARID,
  m_axi_in_18_ARLEN,
  m_axi_in_18_ARLOCK,
  m_axi_in_18_ARPROT,
  m_axi_in_18_ARQOS,
  m_axi_in_18_ARREADY,
  m_axi_in_18_ARSIZE,
  m_axi_in_18_ARVALID,
  m_axi_in_18_AWADDR,
  m_axi_in_18_AWBURST,
  m_axi_in_18_AWCACHE,
  m_axi_in_18_AWID,
  m_axi_in_18_AWLEN,
  m_axi_in_18_AWLOCK,
  m_axi_in_18_AWPROT,
  m_axi_in_18_AWQOS,
  m_axi_in_18_AWREADY,
  m_axi_in_18_AWSIZE,
  m_axi_in_18_AWVALID,
  m_axi_in_18_BID,
  m_axi_in_18_BREADY,
  m_axi_in_18_BRESP,
  m_axi_in_18_BVALID,
  m_axi_in_18_RDATA,
  m_axi_in_18_RID,
  m_axi_in_18_RLAST,
  m_axi_in_18_RREADY,
  m_axi_in_18_RRESP,
  m_axi_in_18_RVALID,
  m_axi_in_18_WDATA,
  m_axi_in_18_WLAST,
  m_axi_in_18_WREADY,
  m_axi_in_18_WSTRB,
  m_axi_in_18_WVALID,
  m_axi_in_19_ARADDR,
  m_axi_in_19_ARBURST,
  m_axi_in_19_ARCACHE,
  m_axi_in_19_ARID,
  m_axi_in_19_ARLEN,
  m_axi_in_19_ARLOCK,
  m_axi_in_19_ARPROT,
  m_axi_in_19_ARQOS,
  m_axi_in_19_ARREADY,
  m_axi_in_19_ARSIZE,
  m_axi_in_19_ARVALID,
  m_axi_in_19_AWADDR,
  m_axi_in_19_AWBURST,
  m_axi_in_19_AWCACHE,
  m_axi_in_19_AWID,
  m_axi_in_19_AWLEN,
  m_axi_in_19_AWLOCK,
  m_axi_in_19_AWPROT,
  m_axi_in_19_AWQOS,
  m_axi_in_19_AWREADY,
  m_axi_in_19_AWSIZE,
  m_axi_in_19_AWVALID,
  m_axi_in_19_BID,
  m_axi_in_19_BREADY,
  m_axi_in_19_BRESP,
  m_axi_in_19_BVALID,
  m_axi_in_19_RDATA,
  m_axi_in_19_RID,
  m_axi_in_19_RLAST,
  m_axi_in_19_RREADY,
  m_axi_in_19_RRESP,
  m_axi_in_19_RVALID,
  m_axi_in_19_WDATA,
  m_axi_in_19_WLAST,
  m_axi_in_19_WREADY,
  m_axi_in_19_WSTRB,
  m_axi_in_19_WVALID,
  m_axi_in_2_ARADDR,
  m_axi_in_2_ARBURST,
  m_axi_in_2_ARCACHE,
  m_axi_in_2_ARID,
  m_axi_in_2_ARLEN,
  m_axi_in_2_ARLOCK,
  m_axi_in_2_ARPROT,
  m_axi_in_2_ARQOS,
  m_axi_in_2_ARREADY,
  m_axi_in_2_ARSIZE,
  m_axi_in_2_ARVALID,
  m_axi_in_2_AWADDR,
  m_axi_in_2_AWBURST,
  m_axi_in_2_AWCACHE,
  m_axi_in_2_AWID,
  m_axi_in_2_AWLEN,
  m_axi_in_2_AWLOCK,
  m_axi_in_2_AWPROT,
  m_axi_in_2_AWQOS,
  m_axi_in_2_AWREADY,
  m_axi_in_2_AWSIZE,
  m_axi_in_2_AWVALID,
  m_axi_in_2_BID,
  m_axi_in_2_BREADY,
  m_axi_in_2_BRESP,
  m_axi_in_2_BVALID,
  m_axi_in_2_RDATA,
  m_axi_in_2_RID,
  m_axi_in_2_RLAST,
  m_axi_in_2_RREADY,
  m_axi_in_2_RRESP,
  m_axi_in_2_RVALID,
  m_axi_in_2_WDATA,
  m_axi_in_2_WLAST,
  m_axi_in_2_WREADY,
  m_axi_in_2_WSTRB,
  m_axi_in_2_WVALID,
  m_axi_in_20_ARADDR,
  m_axi_in_20_ARBURST,
  m_axi_in_20_ARCACHE,
  m_axi_in_20_ARID,
  m_axi_in_20_ARLEN,
  m_axi_in_20_ARLOCK,
  m_axi_in_20_ARPROT,
  m_axi_in_20_ARQOS,
  m_axi_in_20_ARREADY,
  m_axi_in_20_ARSIZE,
  m_axi_in_20_ARVALID,
  m_axi_in_20_AWADDR,
  m_axi_in_20_AWBURST,
  m_axi_in_20_AWCACHE,
  m_axi_in_20_AWID,
  m_axi_in_20_AWLEN,
  m_axi_in_20_AWLOCK,
  m_axi_in_20_AWPROT,
  m_axi_in_20_AWQOS,
  m_axi_in_20_AWREADY,
  m_axi_in_20_AWSIZE,
  m_axi_in_20_AWVALID,
  m_axi_in_20_BID,
  m_axi_in_20_BREADY,
  m_axi_in_20_BRESP,
  m_axi_in_20_BVALID,
  m_axi_in_20_RDATA,
  m_axi_in_20_RID,
  m_axi_in_20_RLAST,
  m_axi_in_20_RREADY,
  m_axi_in_20_RRESP,
  m_axi_in_20_RVALID,
  m_axi_in_20_WDATA,
  m_axi_in_20_WLAST,
  m_axi_in_20_WREADY,
  m_axi_in_20_WSTRB,
  m_axi_in_20_WVALID,
  m_axi_in_21_ARADDR,
  m_axi_in_21_ARBURST,
  m_axi_in_21_ARCACHE,
  m_axi_in_21_ARID,
  m_axi_in_21_ARLEN,
  m_axi_in_21_ARLOCK,
  m_axi_in_21_ARPROT,
  m_axi_in_21_ARQOS,
  m_axi_in_21_ARREADY,
  m_axi_in_21_ARSIZE,
  m_axi_in_21_ARVALID,
  m_axi_in_21_AWADDR,
  m_axi_in_21_AWBURST,
  m_axi_in_21_AWCACHE,
  m_axi_in_21_AWID,
  m_axi_in_21_AWLEN,
  m_axi_in_21_AWLOCK,
  m_axi_in_21_AWPROT,
  m_axi_in_21_AWQOS,
  m_axi_in_21_AWREADY,
  m_axi_in_21_AWSIZE,
  m_axi_in_21_AWVALID,
  m_axi_in_21_BID,
  m_axi_in_21_BREADY,
  m_axi_in_21_BRESP,
  m_axi_in_21_BVALID,
  m_axi_in_21_RDATA,
  m_axi_in_21_RID,
  m_axi_in_21_RLAST,
  m_axi_in_21_RREADY,
  m_axi_in_21_RRESP,
  m_axi_in_21_RVALID,
  m_axi_in_21_WDATA,
  m_axi_in_21_WLAST,
  m_axi_in_21_WREADY,
  m_axi_in_21_WSTRB,
  m_axi_in_21_WVALID,
  m_axi_in_22_ARADDR,
  m_axi_in_22_ARBURST,
  m_axi_in_22_ARCACHE,
  m_axi_in_22_ARID,
  m_axi_in_22_ARLEN,
  m_axi_in_22_ARLOCK,
  m_axi_in_22_ARPROT,
  m_axi_in_22_ARQOS,
  m_axi_in_22_ARREADY,
  m_axi_in_22_ARSIZE,
  m_axi_in_22_ARVALID,
  m_axi_in_22_AWADDR,
  m_axi_in_22_AWBURST,
  m_axi_in_22_AWCACHE,
  m_axi_in_22_AWID,
  m_axi_in_22_AWLEN,
  m_axi_in_22_AWLOCK,
  m_axi_in_22_AWPROT,
  m_axi_in_22_AWQOS,
  m_axi_in_22_AWREADY,
  m_axi_in_22_AWSIZE,
  m_axi_in_22_AWVALID,
  m_axi_in_22_BID,
  m_axi_in_22_BREADY,
  m_axi_in_22_BRESP,
  m_axi_in_22_BVALID,
  m_axi_in_22_RDATA,
  m_axi_in_22_RID,
  m_axi_in_22_RLAST,
  m_axi_in_22_RREADY,
  m_axi_in_22_RRESP,
  m_axi_in_22_RVALID,
  m_axi_in_22_WDATA,
  m_axi_in_22_WLAST,
  m_axi_in_22_WREADY,
  m_axi_in_22_WSTRB,
  m_axi_in_22_WVALID,
  m_axi_in_23_ARADDR,
  m_axi_in_23_ARBURST,
  m_axi_in_23_ARCACHE,
  m_axi_in_23_ARID,
  m_axi_in_23_ARLEN,
  m_axi_in_23_ARLOCK,
  m_axi_in_23_ARPROT,
  m_axi_in_23_ARQOS,
  m_axi_in_23_ARREADY,
  m_axi_in_23_ARSIZE,
  m_axi_in_23_ARVALID,
  m_axi_in_23_AWADDR,
  m_axi_in_23_AWBURST,
  m_axi_in_23_AWCACHE,
  m_axi_in_23_AWID,
  m_axi_in_23_AWLEN,
  m_axi_in_23_AWLOCK,
  m_axi_in_23_AWPROT,
  m_axi_in_23_AWQOS,
  m_axi_in_23_AWREADY,
  m_axi_in_23_AWSIZE,
  m_axi_in_23_AWVALID,
  m_axi_in_23_BID,
  m_axi_in_23_BREADY,
  m_axi_in_23_BRESP,
  m_axi_in_23_BVALID,
  m_axi_in_23_RDATA,
  m_axi_in_23_RID,
  m_axi_in_23_RLAST,
  m_axi_in_23_RREADY,
  m_axi_in_23_RRESP,
  m_axi_in_23_RVALID,
  m_axi_in_23_WDATA,
  m_axi_in_23_WLAST,
  m_axi_in_23_WREADY,
  m_axi_in_23_WSTRB,
  m_axi_in_23_WVALID,
  m_axi_in_24_ARADDR,
  m_axi_in_24_ARBURST,
  m_axi_in_24_ARCACHE,
  m_axi_in_24_ARID,
  m_axi_in_24_ARLEN,
  m_axi_in_24_ARLOCK,
  m_axi_in_24_ARPROT,
  m_axi_in_24_ARQOS,
  m_axi_in_24_ARREADY,
  m_axi_in_24_ARSIZE,
  m_axi_in_24_ARVALID,
  m_axi_in_24_AWADDR,
  m_axi_in_24_AWBURST,
  m_axi_in_24_AWCACHE,
  m_axi_in_24_AWID,
  m_axi_in_24_AWLEN,
  m_axi_in_24_AWLOCK,
  m_axi_in_24_AWPROT,
  m_axi_in_24_AWQOS,
  m_axi_in_24_AWREADY,
  m_axi_in_24_AWSIZE,
  m_axi_in_24_AWVALID,
  m_axi_in_24_BID,
  m_axi_in_24_BREADY,
  m_axi_in_24_BRESP,
  m_axi_in_24_BVALID,
  m_axi_in_24_RDATA,
  m_axi_in_24_RID,
  m_axi_in_24_RLAST,
  m_axi_in_24_RREADY,
  m_axi_in_24_RRESP,
  m_axi_in_24_RVALID,
  m_axi_in_24_WDATA,
  m_axi_in_24_WLAST,
  m_axi_in_24_WREADY,
  m_axi_in_24_WSTRB,
  m_axi_in_24_WVALID,
  m_axi_in_25_ARADDR,
  m_axi_in_25_ARBURST,
  m_axi_in_25_ARCACHE,
  m_axi_in_25_ARID,
  m_axi_in_25_ARLEN,
  m_axi_in_25_ARLOCK,
  m_axi_in_25_ARPROT,
  m_axi_in_25_ARQOS,
  m_axi_in_25_ARREADY,
  m_axi_in_25_ARSIZE,
  m_axi_in_25_ARVALID,
  m_axi_in_25_AWADDR,
  m_axi_in_25_AWBURST,
  m_axi_in_25_AWCACHE,
  m_axi_in_25_AWID,
  m_axi_in_25_AWLEN,
  m_axi_in_25_AWLOCK,
  m_axi_in_25_AWPROT,
  m_axi_in_25_AWQOS,
  m_axi_in_25_AWREADY,
  m_axi_in_25_AWSIZE,
  m_axi_in_25_AWVALID,
  m_axi_in_25_BID,
  m_axi_in_25_BREADY,
  m_axi_in_25_BRESP,
  m_axi_in_25_BVALID,
  m_axi_in_25_RDATA,
  m_axi_in_25_RID,
  m_axi_in_25_RLAST,
  m_axi_in_25_RREADY,
  m_axi_in_25_RRESP,
  m_axi_in_25_RVALID,
  m_axi_in_25_WDATA,
  m_axi_in_25_WLAST,
  m_axi_in_25_WREADY,
  m_axi_in_25_WSTRB,
  m_axi_in_25_WVALID,
  m_axi_in_26_ARADDR,
  m_axi_in_26_ARBURST,
  m_axi_in_26_ARCACHE,
  m_axi_in_26_ARID,
  m_axi_in_26_ARLEN,
  m_axi_in_26_ARLOCK,
  m_axi_in_26_ARPROT,
  m_axi_in_26_ARQOS,
  m_axi_in_26_ARREADY,
  m_axi_in_26_ARSIZE,
  m_axi_in_26_ARVALID,
  m_axi_in_26_AWADDR,
  m_axi_in_26_AWBURST,
  m_axi_in_26_AWCACHE,
  m_axi_in_26_AWID,
  m_axi_in_26_AWLEN,
  m_axi_in_26_AWLOCK,
  m_axi_in_26_AWPROT,
  m_axi_in_26_AWQOS,
  m_axi_in_26_AWREADY,
  m_axi_in_26_AWSIZE,
  m_axi_in_26_AWVALID,
  m_axi_in_26_BID,
  m_axi_in_26_BREADY,
  m_axi_in_26_BRESP,
  m_axi_in_26_BVALID,
  m_axi_in_26_RDATA,
  m_axi_in_26_RID,
  m_axi_in_26_RLAST,
  m_axi_in_26_RREADY,
  m_axi_in_26_RRESP,
  m_axi_in_26_RVALID,
  m_axi_in_26_WDATA,
  m_axi_in_26_WLAST,
  m_axi_in_26_WREADY,
  m_axi_in_26_WSTRB,
  m_axi_in_26_WVALID,
  m_axi_in_27_ARADDR,
  m_axi_in_27_ARBURST,
  m_axi_in_27_ARCACHE,
  m_axi_in_27_ARID,
  m_axi_in_27_ARLEN,
  m_axi_in_27_ARLOCK,
  m_axi_in_27_ARPROT,
  m_axi_in_27_ARQOS,
  m_axi_in_27_ARREADY,
  m_axi_in_27_ARSIZE,
  m_axi_in_27_ARVALID,
  m_axi_in_27_AWADDR,
  m_axi_in_27_AWBURST,
  m_axi_in_27_AWCACHE,
  m_axi_in_27_AWID,
  m_axi_in_27_AWLEN,
  m_axi_in_27_AWLOCK,
  m_axi_in_27_AWPROT,
  m_axi_in_27_AWQOS,
  m_axi_in_27_AWREADY,
  m_axi_in_27_AWSIZE,
  m_axi_in_27_AWVALID,
  m_axi_in_27_BID,
  m_axi_in_27_BREADY,
  m_axi_in_27_BRESP,
  m_axi_in_27_BVALID,
  m_axi_in_27_RDATA,
  m_axi_in_27_RID,
  m_axi_in_27_RLAST,
  m_axi_in_27_RREADY,
  m_axi_in_27_RRESP,
  m_axi_in_27_RVALID,
  m_axi_in_27_WDATA,
  m_axi_in_27_WLAST,
  m_axi_in_27_WREADY,
  m_axi_in_27_WSTRB,
  m_axi_in_27_WVALID,
  m_axi_in_28_ARADDR,
  m_axi_in_28_ARBURST,
  m_axi_in_28_ARCACHE,
  m_axi_in_28_ARID,
  m_axi_in_28_ARLEN,
  m_axi_in_28_ARLOCK,
  m_axi_in_28_ARPROT,
  m_axi_in_28_ARQOS,
  m_axi_in_28_ARREADY,
  m_axi_in_28_ARSIZE,
  m_axi_in_28_ARVALID,
  m_axi_in_28_AWADDR,
  m_axi_in_28_AWBURST,
  m_axi_in_28_AWCACHE,
  m_axi_in_28_AWID,
  m_axi_in_28_AWLEN,
  m_axi_in_28_AWLOCK,
  m_axi_in_28_AWPROT,
  m_axi_in_28_AWQOS,
  m_axi_in_28_AWREADY,
  m_axi_in_28_AWSIZE,
  m_axi_in_28_AWVALID,
  m_axi_in_28_BID,
  m_axi_in_28_BREADY,
  m_axi_in_28_BRESP,
  m_axi_in_28_BVALID,
  m_axi_in_28_RDATA,
  m_axi_in_28_RID,
  m_axi_in_28_RLAST,
  m_axi_in_28_RREADY,
  m_axi_in_28_RRESP,
  m_axi_in_28_RVALID,
  m_axi_in_28_WDATA,
  m_axi_in_28_WLAST,
  m_axi_in_28_WREADY,
  m_axi_in_28_WSTRB,
  m_axi_in_28_WVALID,
  m_axi_in_29_ARADDR,
  m_axi_in_29_ARBURST,
  m_axi_in_29_ARCACHE,
  m_axi_in_29_ARID,
  m_axi_in_29_ARLEN,
  m_axi_in_29_ARLOCK,
  m_axi_in_29_ARPROT,
  m_axi_in_29_ARQOS,
  m_axi_in_29_ARREADY,
  m_axi_in_29_ARSIZE,
  m_axi_in_29_ARVALID,
  m_axi_in_29_AWADDR,
  m_axi_in_29_AWBURST,
  m_axi_in_29_AWCACHE,
  m_axi_in_29_AWID,
  m_axi_in_29_AWLEN,
  m_axi_in_29_AWLOCK,
  m_axi_in_29_AWPROT,
  m_axi_in_29_AWQOS,
  m_axi_in_29_AWREADY,
  m_axi_in_29_AWSIZE,
  m_axi_in_29_AWVALID,
  m_axi_in_29_BID,
  m_axi_in_29_BREADY,
  m_axi_in_29_BRESP,
  m_axi_in_29_BVALID,
  m_axi_in_29_RDATA,
  m_axi_in_29_RID,
  m_axi_in_29_RLAST,
  m_axi_in_29_RREADY,
  m_axi_in_29_RRESP,
  m_axi_in_29_RVALID,
  m_axi_in_29_WDATA,
  m_axi_in_29_WLAST,
  m_axi_in_29_WREADY,
  m_axi_in_29_WSTRB,
  m_axi_in_29_WVALID,
  m_axi_in_3_ARADDR,
  m_axi_in_3_ARBURST,
  m_axi_in_3_ARCACHE,
  m_axi_in_3_ARID,
  m_axi_in_3_ARLEN,
  m_axi_in_3_ARLOCK,
  m_axi_in_3_ARPROT,
  m_axi_in_3_ARQOS,
  m_axi_in_3_ARREADY,
  m_axi_in_3_ARSIZE,
  m_axi_in_3_ARVALID,
  m_axi_in_3_AWADDR,
  m_axi_in_3_AWBURST,
  m_axi_in_3_AWCACHE,
  m_axi_in_3_AWID,
  m_axi_in_3_AWLEN,
  m_axi_in_3_AWLOCK,
  m_axi_in_3_AWPROT,
  m_axi_in_3_AWQOS,
  m_axi_in_3_AWREADY,
  m_axi_in_3_AWSIZE,
  m_axi_in_3_AWVALID,
  m_axi_in_3_BID,
  m_axi_in_3_BREADY,
  m_axi_in_3_BRESP,
  m_axi_in_3_BVALID,
  m_axi_in_3_RDATA,
  m_axi_in_3_RID,
  m_axi_in_3_RLAST,
  m_axi_in_3_RREADY,
  m_axi_in_3_RRESP,
  m_axi_in_3_RVALID,
  m_axi_in_3_WDATA,
  m_axi_in_3_WLAST,
  m_axi_in_3_WREADY,
  m_axi_in_3_WSTRB,
  m_axi_in_3_WVALID,
  m_axi_in_30_ARADDR,
  m_axi_in_30_ARBURST,
  m_axi_in_30_ARCACHE,
  m_axi_in_30_ARID,
  m_axi_in_30_ARLEN,
  m_axi_in_30_ARLOCK,
  m_axi_in_30_ARPROT,
  m_axi_in_30_ARQOS,
  m_axi_in_30_ARREADY,
  m_axi_in_30_ARSIZE,
  m_axi_in_30_ARVALID,
  m_axi_in_30_AWADDR,
  m_axi_in_30_AWBURST,
  m_axi_in_30_AWCACHE,
  m_axi_in_30_AWID,
  m_axi_in_30_AWLEN,
  m_axi_in_30_AWLOCK,
  m_axi_in_30_AWPROT,
  m_axi_in_30_AWQOS,
  m_axi_in_30_AWREADY,
  m_axi_in_30_AWSIZE,
  m_axi_in_30_AWVALID,
  m_axi_in_30_BID,
  m_axi_in_30_BREADY,
  m_axi_in_30_BRESP,
  m_axi_in_30_BVALID,
  m_axi_in_30_RDATA,
  m_axi_in_30_RID,
  m_axi_in_30_RLAST,
  m_axi_in_30_RREADY,
  m_axi_in_30_RRESP,
  m_axi_in_30_RVALID,
  m_axi_in_30_WDATA,
  m_axi_in_30_WLAST,
  m_axi_in_30_WREADY,
  m_axi_in_30_WSTRB,
  m_axi_in_30_WVALID,
  m_axi_in_31_ARADDR,
  m_axi_in_31_ARBURST,
  m_axi_in_31_ARCACHE,
  m_axi_in_31_ARID,
  m_axi_in_31_ARLEN,
  m_axi_in_31_ARLOCK,
  m_axi_in_31_ARPROT,
  m_axi_in_31_ARQOS,
  m_axi_in_31_ARREADY,
  m_axi_in_31_ARSIZE,
  m_axi_in_31_ARVALID,
  m_axi_in_31_AWADDR,
  m_axi_in_31_AWBURST,
  m_axi_in_31_AWCACHE,
  m_axi_in_31_AWID,
  m_axi_in_31_AWLEN,
  m_axi_in_31_AWLOCK,
  m_axi_in_31_AWPROT,
  m_axi_in_31_AWQOS,
  m_axi_in_31_AWREADY,
  m_axi_in_31_AWSIZE,
  m_axi_in_31_AWVALID,
  m_axi_in_31_BID,
  m_axi_in_31_BREADY,
  m_axi_in_31_BRESP,
  m_axi_in_31_BVALID,
  m_axi_in_31_RDATA,
  m_axi_in_31_RID,
  m_axi_in_31_RLAST,
  m_axi_in_31_RREADY,
  m_axi_in_31_RRESP,
  m_axi_in_31_RVALID,
  m_axi_in_31_WDATA,
  m_axi_in_31_WLAST,
  m_axi_in_31_WREADY,
  m_axi_in_31_WSTRB,
  m_axi_in_31_WVALID,
  m_axi_in_32_ARADDR,
  m_axi_in_32_ARBURST,
  m_axi_in_32_ARCACHE,
  m_axi_in_32_ARID,
  m_axi_in_32_ARLEN,
  m_axi_in_32_ARLOCK,
  m_axi_in_32_ARPROT,
  m_axi_in_32_ARQOS,
  m_axi_in_32_ARREADY,
  m_axi_in_32_ARSIZE,
  m_axi_in_32_ARVALID,
  m_axi_in_32_AWADDR,
  m_axi_in_32_AWBURST,
  m_axi_in_32_AWCACHE,
  m_axi_in_32_AWID,
  m_axi_in_32_AWLEN,
  m_axi_in_32_AWLOCK,
  m_axi_in_32_AWPROT,
  m_axi_in_32_AWQOS,
  m_axi_in_32_AWREADY,
  m_axi_in_32_AWSIZE,
  m_axi_in_32_AWVALID,
  m_axi_in_32_BID,
  m_axi_in_32_BREADY,
  m_axi_in_32_BRESP,
  m_axi_in_32_BVALID,
  m_axi_in_32_RDATA,
  m_axi_in_32_RID,
  m_axi_in_32_RLAST,
  m_axi_in_32_RREADY,
  m_axi_in_32_RRESP,
  m_axi_in_32_RVALID,
  m_axi_in_32_WDATA,
  m_axi_in_32_WLAST,
  m_axi_in_32_WREADY,
  m_axi_in_32_WSTRB,
  m_axi_in_32_WVALID,
  m_axi_in_33_ARADDR,
  m_axi_in_33_ARBURST,
  m_axi_in_33_ARCACHE,
  m_axi_in_33_ARID,
  m_axi_in_33_ARLEN,
  m_axi_in_33_ARLOCK,
  m_axi_in_33_ARPROT,
  m_axi_in_33_ARQOS,
  m_axi_in_33_ARREADY,
  m_axi_in_33_ARSIZE,
  m_axi_in_33_ARVALID,
  m_axi_in_33_AWADDR,
  m_axi_in_33_AWBURST,
  m_axi_in_33_AWCACHE,
  m_axi_in_33_AWID,
  m_axi_in_33_AWLEN,
  m_axi_in_33_AWLOCK,
  m_axi_in_33_AWPROT,
  m_axi_in_33_AWQOS,
  m_axi_in_33_AWREADY,
  m_axi_in_33_AWSIZE,
  m_axi_in_33_AWVALID,
  m_axi_in_33_BID,
  m_axi_in_33_BREADY,
  m_axi_in_33_BRESP,
  m_axi_in_33_BVALID,
  m_axi_in_33_RDATA,
  m_axi_in_33_RID,
  m_axi_in_33_RLAST,
  m_axi_in_33_RREADY,
  m_axi_in_33_RRESP,
  m_axi_in_33_RVALID,
  m_axi_in_33_WDATA,
  m_axi_in_33_WLAST,
  m_axi_in_33_WREADY,
  m_axi_in_33_WSTRB,
  m_axi_in_33_WVALID,
  m_axi_in_34_ARADDR,
  m_axi_in_34_ARBURST,
  m_axi_in_34_ARCACHE,
  m_axi_in_34_ARID,
  m_axi_in_34_ARLEN,
  m_axi_in_34_ARLOCK,
  m_axi_in_34_ARPROT,
  m_axi_in_34_ARQOS,
  m_axi_in_34_ARREADY,
  m_axi_in_34_ARSIZE,
  m_axi_in_34_ARVALID,
  m_axi_in_34_AWADDR,
  m_axi_in_34_AWBURST,
  m_axi_in_34_AWCACHE,
  m_axi_in_34_AWID,
  m_axi_in_34_AWLEN,
  m_axi_in_34_AWLOCK,
  m_axi_in_34_AWPROT,
  m_axi_in_34_AWQOS,
  m_axi_in_34_AWREADY,
  m_axi_in_34_AWSIZE,
  m_axi_in_34_AWVALID,
  m_axi_in_34_BID,
  m_axi_in_34_BREADY,
  m_axi_in_34_BRESP,
  m_axi_in_34_BVALID,
  m_axi_in_34_RDATA,
  m_axi_in_34_RID,
  m_axi_in_34_RLAST,
  m_axi_in_34_RREADY,
  m_axi_in_34_RRESP,
  m_axi_in_34_RVALID,
  m_axi_in_34_WDATA,
  m_axi_in_34_WLAST,
  m_axi_in_34_WREADY,
  m_axi_in_34_WSTRB,
  m_axi_in_34_WVALID,
  m_axi_in_35_ARADDR,
  m_axi_in_35_ARBURST,
  m_axi_in_35_ARCACHE,
  m_axi_in_35_ARID,
  m_axi_in_35_ARLEN,
  m_axi_in_35_ARLOCK,
  m_axi_in_35_ARPROT,
  m_axi_in_35_ARQOS,
  m_axi_in_35_ARREADY,
  m_axi_in_35_ARSIZE,
  m_axi_in_35_ARVALID,
  m_axi_in_35_AWADDR,
  m_axi_in_35_AWBURST,
  m_axi_in_35_AWCACHE,
  m_axi_in_35_AWID,
  m_axi_in_35_AWLEN,
  m_axi_in_35_AWLOCK,
  m_axi_in_35_AWPROT,
  m_axi_in_35_AWQOS,
  m_axi_in_35_AWREADY,
  m_axi_in_35_AWSIZE,
  m_axi_in_35_AWVALID,
  m_axi_in_35_BID,
  m_axi_in_35_BREADY,
  m_axi_in_35_BRESP,
  m_axi_in_35_BVALID,
  m_axi_in_35_RDATA,
  m_axi_in_35_RID,
  m_axi_in_35_RLAST,
  m_axi_in_35_RREADY,
  m_axi_in_35_RRESP,
  m_axi_in_35_RVALID,
  m_axi_in_35_WDATA,
  m_axi_in_35_WLAST,
  m_axi_in_35_WREADY,
  m_axi_in_35_WSTRB,
  m_axi_in_35_WVALID,
  m_axi_in_36_ARADDR,
  m_axi_in_36_ARBURST,
  m_axi_in_36_ARCACHE,
  m_axi_in_36_ARID,
  m_axi_in_36_ARLEN,
  m_axi_in_36_ARLOCK,
  m_axi_in_36_ARPROT,
  m_axi_in_36_ARQOS,
  m_axi_in_36_ARREADY,
  m_axi_in_36_ARSIZE,
  m_axi_in_36_ARVALID,
  m_axi_in_36_AWADDR,
  m_axi_in_36_AWBURST,
  m_axi_in_36_AWCACHE,
  m_axi_in_36_AWID,
  m_axi_in_36_AWLEN,
  m_axi_in_36_AWLOCK,
  m_axi_in_36_AWPROT,
  m_axi_in_36_AWQOS,
  m_axi_in_36_AWREADY,
  m_axi_in_36_AWSIZE,
  m_axi_in_36_AWVALID,
  m_axi_in_36_BID,
  m_axi_in_36_BREADY,
  m_axi_in_36_BRESP,
  m_axi_in_36_BVALID,
  m_axi_in_36_RDATA,
  m_axi_in_36_RID,
  m_axi_in_36_RLAST,
  m_axi_in_36_RREADY,
  m_axi_in_36_RRESP,
  m_axi_in_36_RVALID,
  m_axi_in_36_WDATA,
  m_axi_in_36_WLAST,
  m_axi_in_36_WREADY,
  m_axi_in_36_WSTRB,
  m_axi_in_36_WVALID,
  m_axi_in_37_ARADDR,
  m_axi_in_37_ARBURST,
  m_axi_in_37_ARCACHE,
  m_axi_in_37_ARID,
  m_axi_in_37_ARLEN,
  m_axi_in_37_ARLOCK,
  m_axi_in_37_ARPROT,
  m_axi_in_37_ARQOS,
  m_axi_in_37_ARREADY,
  m_axi_in_37_ARSIZE,
  m_axi_in_37_ARVALID,
  m_axi_in_37_AWADDR,
  m_axi_in_37_AWBURST,
  m_axi_in_37_AWCACHE,
  m_axi_in_37_AWID,
  m_axi_in_37_AWLEN,
  m_axi_in_37_AWLOCK,
  m_axi_in_37_AWPROT,
  m_axi_in_37_AWQOS,
  m_axi_in_37_AWREADY,
  m_axi_in_37_AWSIZE,
  m_axi_in_37_AWVALID,
  m_axi_in_37_BID,
  m_axi_in_37_BREADY,
  m_axi_in_37_BRESP,
  m_axi_in_37_BVALID,
  m_axi_in_37_RDATA,
  m_axi_in_37_RID,
  m_axi_in_37_RLAST,
  m_axi_in_37_RREADY,
  m_axi_in_37_RRESP,
  m_axi_in_37_RVALID,
  m_axi_in_37_WDATA,
  m_axi_in_37_WLAST,
  m_axi_in_37_WREADY,
  m_axi_in_37_WSTRB,
  m_axi_in_37_WVALID,
  m_axi_in_38_ARADDR,
  m_axi_in_38_ARBURST,
  m_axi_in_38_ARCACHE,
  m_axi_in_38_ARID,
  m_axi_in_38_ARLEN,
  m_axi_in_38_ARLOCK,
  m_axi_in_38_ARPROT,
  m_axi_in_38_ARQOS,
  m_axi_in_38_ARREADY,
  m_axi_in_38_ARSIZE,
  m_axi_in_38_ARVALID,
  m_axi_in_38_AWADDR,
  m_axi_in_38_AWBURST,
  m_axi_in_38_AWCACHE,
  m_axi_in_38_AWID,
  m_axi_in_38_AWLEN,
  m_axi_in_38_AWLOCK,
  m_axi_in_38_AWPROT,
  m_axi_in_38_AWQOS,
  m_axi_in_38_AWREADY,
  m_axi_in_38_AWSIZE,
  m_axi_in_38_AWVALID,
  m_axi_in_38_BID,
  m_axi_in_38_BREADY,
  m_axi_in_38_BRESP,
  m_axi_in_38_BVALID,
  m_axi_in_38_RDATA,
  m_axi_in_38_RID,
  m_axi_in_38_RLAST,
  m_axi_in_38_RREADY,
  m_axi_in_38_RRESP,
  m_axi_in_38_RVALID,
  m_axi_in_38_WDATA,
  m_axi_in_38_WLAST,
  m_axi_in_38_WREADY,
  m_axi_in_38_WSTRB,
  m_axi_in_38_WVALID,
  m_axi_in_39_ARADDR,
  m_axi_in_39_ARBURST,
  m_axi_in_39_ARCACHE,
  m_axi_in_39_ARID,
  m_axi_in_39_ARLEN,
  m_axi_in_39_ARLOCK,
  m_axi_in_39_ARPROT,
  m_axi_in_39_ARQOS,
  m_axi_in_39_ARREADY,
  m_axi_in_39_ARSIZE,
  m_axi_in_39_ARVALID,
  m_axi_in_39_AWADDR,
  m_axi_in_39_AWBURST,
  m_axi_in_39_AWCACHE,
  m_axi_in_39_AWID,
  m_axi_in_39_AWLEN,
  m_axi_in_39_AWLOCK,
  m_axi_in_39_AWPROT,
  m_axi_in_39_AWQOS,
  m_axi_in_39_AWREADY,
  m_axi_in_39_AWSIZE,
  m_axi_in_39_AWVALID,
  m_axi_in_39_BID,
  m_axi_in_39_BREADY,
  m_axi_in_39_BRESP,
  m_axi_in_39_BVALID,
  m_axi_in_39_RDATA,
  m_axi_in_39_RID,
  m_axi_in_39_RLAST,
  m_axi_in_39_RREADY,
  m_axi_in_39_RRESP,
  m_axi_in_39_RVALID,
  m_axi_in_39_WDATA,
  m_axi_in_39_WLAST,
  m_axi_in_39_WREADY,
  m_axi_in_39_WSTRB,
  m_axi_in_39_WVALID,
  m_axi_in_4_ARADDR,
  m_axi_in_4_ARBURST,
  m_axi_in_4_ARCACHE,
  m_axi_in_4_ARID,
  m_axi_in_4_ARLEN,
  m_axi_in_4_ARLOCK,
  m_axi_in_4_ARPROT,
  m_axi_in_4_ARQOS,
  m_axi_in_4_ARREADY,
  m_axi_in_4_ARSIZE,
  m_axi_in_4_ARVALID,
  m_axi_in_4_AWADDR,
  m_axi_in_4_AWBURST,
  m_axi_in_4_AWCACHE,
  m_axi_in_4_AWID,
  m_axi_in_4_AWLEN,
  m_axi_in_4_AWLOCK,
  m_axi_in_4_AWPROT,
  m_axi_in_4_AWQOS,
  m_axi_in_4_AWREADY,
  m_axi_in_4_AWSIZE,
  m_axi_in_4_AWVALID,
  m_axi_in_4_BID,
  m_axi_in_4_BREADY,
  m_axi_in_4_BRESP,
  m_axi_in_4_BVALID,
  m_axi_in_4_RDATA,
  m_axi_in_4_RID,
  m_axi_in_4_RLAST,
  m_axi_in_4_RREADY,
  m_axi_in_4_RRESP,
  m_axi_in_4_RVALID,
  m_axi_in_4_WDATA,
  m_axi_in_4_WLAST,
  m_axi_in_4_WREADY,
  m_axi_in_4_WSTRB,
  m_axi_in_4_WVALID,
  m_axi_in_40_ARADDR,
  m_axi_in_40_ARBURST,
  m_axi_in_40_ARCACHE,
  m_axi_in_40_ARID,
  m_axi_in_40_ARLEN,
  m_axi_in_40_ARLOCK,
  m_axi_in_40_ARPROT,
  m_axi_in_40_ARQOS,
  m_axi_in_40_ARREADY,
  m_axi_in_40_ARSIZE,
  m_axi_in_40_ARVALID,
  m_axi_in_40_AWADDR,
  m_axi_in_40_AWBURST,
  m_axi_in_40_AWCACHE,
  m_axi_in_40_AWID,
  m_axi_in_40_AWLEN,
  m_axi_in_40_AWLOCK,
  m_axi_in_40_AWPROT,
  m_axi_in_40_AWQOS,
  m_axi_in_40_AWREADY,
  m_axi_in_40_AWSIZE,
  m_axi_in_40_AWVALID,
  m_axi_in_40_BID,
  m_axi_in_40_BREADY,
  m_axi_in_40_BRESP,
  m_axi_in_40_BVALID,
  m_axi_in_40_RDATA,
  m_axi_in_40_RID,
  m_axi_in_40_RLAST,
  m_axi_in_40_RREADY,
  m_axi_in_40_RRESP,
  m_axi_in_40_RVALID,
  m_axi_in_40_WDATA,
  m_axi_in_40_WLAST,
  m_axi_in_40_WREADY,
  m_axi_in_40_WSTRB,
  m_axi_in_40_WVALID,
  m_axi_in_41_ARADDR,
  m_axi_in_41_ARBURST,
  m_axi_in_41_ARCACHE,
  m_axi_in_41_ARID,
  m_axi_in_41_ARLEN,
  m_axi_in_41_ARLOCK,
  m_axi_in_41_ARPROT,
  m_axi_in_41_ARQOS,
  m_axi_in_41_ARREADY,
  m_axi_in_41_ARSIZE,
  m_axi_in_41_ARVALID,
  m_axi_in_41_AWADDR,
  m_axi_in_41_AWBURST,
  m_axi_in_41_AWCACHE,
  m_axi_in_41_AWID,
  m_axi_in_41_AWLEN,
  m_axi_in_41_AWLOCK,
  m_axi_in_41_AWPROT,
  m_axi_in_41_AWQOS,
  m_axi_in_41_AWREADY,
  m_axi_in_41_AWSIZE,
  m_axi_in_41_AWVALID,
  m_axi_in_41_BID,
  m_axi_in_41_BREADY,
  m_axi_in_41_BRESP,
  m_axi_in_41_BVALID,
  m_axi_in_41_RDATA,
  m_axi_in_41_RID,
  m_axi_in_41_RLAST,
  m_axi_in_41_RREADY,
  m_axi_in_41_RRESP,
  m_axi_in_41_RVALID,
  m_axi_in_41_WDATA,
  m_axi_in_41_WLAST,
  m_axi_in_41_WREADY,
  m_axi_in_41_WSTRB,
  m_axi_in_41_WVALID,
  m_axi_in_42_ARADDR,
  m_axi_in_42_ARBURST,
  m_axi_in_42_ARCACHE,
  m_axi_in_42_ARID,
  m_axi_in_42_ARLEN,
  m_axi_in_42_ARLOCK,
  m_axi_in_42_ARPROT,
  m_axi_in_42_ARQOS,
  m_axi_in_42_ARREADY,
  m_axi_in_42_ARSIZE,
  m_axi_in_42_ARVALID,
  m_axi_in_42_AWADDR,
  m_axi_in_42_AWBURST,
  m_axi_in_42_AWCACHE,
  m_axi_in_42_AWID,
  m_axi_in_42_AWLEN,
  m_axi_in_42_AWLOCK,
  m_axi_in_42_AWPROT,
  m_axi_in_42_AWQOS,
  m_axi_in_42_AWREADY,
  m_axi_in_42_AWSIZE,
  m_axi_in_42_AWVALID,
  m_axi_in_42_BID,
  m_axi_in_42_BREADY,
  m_axi_in_42_BRESP,
  m_axi_in_42_BVALID,
  m_axi_in_42_RDATA,
  m_axi_in_42_RID,
  m_axi_in_42_RLAST,
  m_axi_in_42_RREADY,
  m_axi_in_42_RRESP,
  m_axi_in_42_RVALID,
  m_axi_in_42_WDATA,
  m_axi_in_42_WLAST,
  m_axi_in_42_WREADY,
  m_axi_in_42_WSTRB,
  m_axi_in_42_WVALID,
  m_axi_in_43_ARADDR,
  m_axi_in_43_ARBURST,
  m_axi_in_43_ARCACHE,
  m_axi_in_43_ARID,
  m_axi_in_43_ARLEN,
  m_axi_in_43_ARLOCK,
  m_axi_in_43_ARPROT,
  m_axi_in_43_ARQOS,
  m_axi_in_43_ARREADY,
  m_axi_in_43_ARSIZE,
  m_axi_in_43_ARVALID,
  m_axi_in_43_AWADDR,
  m_axi_in_43_AWBURST,
  m_axi_in_43_AWCACHE,
  m_axi_in_43_AWID,
  m_axi_in_43_AWLEN,
  m_axi_in_43_AWLOCK,
  m_axi_in_43_AWPROT,
  m_axi_in_43_AWQOS,
  m_axi_in_43_AWREADY,
  m_axi_in_43_AWSIZE,
  m_axi_in_43_AWVALID,
  m_axi_in_43_BID,
  m_axi_in_43_BREADY,
  m_axi_in_43_BRESP,
  m_axi_in_43_BVALID,
  m_axi_in_43_RDATA,
  m_axi_in_43_RID,
  m_axi_in_43_RLAST,
  m_axi_in_43_RREADY,
  m_axi_in_43_RRESP,
  m_axi_in_43_RVALID,
  m_axi_in_43_WDATA,
  m_axi_in_43_WLAST,
  m_axi_in_43_WREADY,
  m_axi_in_43_WSTRB,
  m_axi_in_43_WVALID,
  m_axi_in_44_ARADDR,
  m_axi_in_44_ARBURST,
  m_axi_in_44_ARCACHE,
  m_axi_in_44_ARID,
  m_axi_in_44_ARLEN,
  m_axi_in_44_ARLOCK,
  m_axi_in_44_ARPROT,
  m_axi_in_44_ARQOS,
  m_axi_in_44_ARREADY,
  m_axi_in_44_ARSIZE,
  m_axi_in_44_ARVALID,
  m_axi_in_44_AWADDR,
  m_axi_in_44_AWBURST,
  m_axi_in_44_AWCACHE,
  m_axi_in_44_AWID,
  m_axi_in_44_AWLEN,
  m_axi_in_44_AWLOCK,
  m_axi_in_44_AWPROT,
  m_axi_in_44_AWQOS,
  m_axi_in_44_AWREADY,
  m_axi_in_44_AWSIZE,
  m_axi_in_44_AWVALID,
  m_axi_in_44_BID,
  m_axi_in_44_BREADY,
  m_axi_in_44_BRESP,
  m_axi_in_44_BVALID,
  m_axi_in_44_RDATA,
  m_axi_in_44_RID,
  m_axi_in_44_RLAST,
  m_axi_in_44_RREADY,
  m_axi_in_44_RRESP,
  m_axi_in_44_RVALID,
  m_axi_in_44_WDATA,
  m_axi_in_44_WLAST,
  m_axi_in_44_WREADY,
  m_axi_in_44_WSTRB,
  m_axi_in_44_WVALID,
  m_axi_in_45_ARADDR,
  m_axi_in_45_ARBURST,
  m_axi_in_45_ARCACHE,
  m_axi_in_45_ARID,
  m_axi_in_45_ARLEN,
  m_axi_in_45_ARLOCK,
  m_axi_in_45_ARPROT,
  m_axi_in_45_ARQOS,
  m_axi_in_45_ARREADY,
  m_axi_in_45_ARSIZE,
  m_axi_in_45_ARVALID,
  m_axi_in_45_AWADDR,
  m_axi_in_45_AWBURST,
  m_axi_in_45_AWCACHE,
  m_axi_in_45_AWID,
  m_axi_in_45_AWLEN,
  m_axi_in_45_AWLOCK,
  m_axi_in_45_AWPROT,
  m_axi_in_45_AWQOS,
  m_axi_in_45_AWREADY,
  m_axi_in_45_AWSIZE,
  m_axi_in_45_AWVALID,
  m_axi_in_45_BID,
  m_axi_in_45_BREADY,
  m_axi_in_45_BRESP,
  m_axi_in_45_BVALID,
  m_axi_in_45_RDATA,
  m_axi_in_45_RID,
  m_axi_in_45_RLAST,
  m_axi_in_45_RREADY,
  m_axi_in_45_RRESP,
  m_axi_in_45_RVALID,
  m_axi_in_45_WDATA,
  m_axi_in_45_WLAST,
  m_axi_in_45_WREADY,
  m_axi_in_45_WSTRB,
  m_axi_in_45_WVALID,
  m_axi_in_46_ARADDR,
  m_axi_in_46_ARBURST,
  m_axi_in_46_ARCACHE,
  m_axi_in_46_ARID,
  m_axi_in_46_ARLEN,
  m_axi_in_46_ARLOCK,
  m_axi_in_46_ARPROT,
  m_axi_in_46_ARQOS,
  m_axi_in_46_ARREADY,
  m_axi_in_46_ARSIZE,
  m_axi_in_46_ARVALID,
  m_axi_in_46_AWADDR,
  m_axi_in_46_AWBURST,
  m_axi_in_46_AWCACHE,
  m_axi_in_46_AWID,
  m_axi_in_46_AWLEN,
  m_axi_in_46_AWLOCK,
  m_axi_in_46_AWPROT,
  m_axi_in_46_AWQOS,
  m_axi_in_46_AWREADY,
  m_axi_in_46_AWSIZE,
  m_axi_in_46_AWVALID,
  m_axi_in_46_BID,
  m_axi_in_46_BREADY,
  m_axi_in_46_BRESP,
  m_axi_in_46_BVALID,
  m_axi_in_46_RDATA,
  m_axi_in_46_RID,
  m_axi_in_46_RLAST,
  m_axi_in_46_RREADY,
  m_axi_in_46_RRESP,
  m_axi_in_46_RVALID,
  m_axi_in_46_WDATA,
  m_axi_in_46_WLAST,
  m_axi_in_46_WREADY,
  m_axi_in_46_WSTRB,
  m_axi_in_46_WVALID,
  m_axi_in_47_ARADDR,
  m_axi_in_47_ARBURST,
  m_axi_in_47_ARCACHE,
  m_axi_in_47_ARID,
  m_axi_in_47_ARLEN,
  m_axi_in_47_ARLOCK,
  m_axi_in_47_ARPROT,
  m_axi_in_47_ARQOS,
  m_axi_in_47_ARREADY,
  m_axi_in_47_ARSIZE,
  m_axi_in_47_ARVALID,
  m_axi_in_47_AWADDR,
  m_axi_in_47_AWBURST,
  m_axi_in_47_AWCACHE,
  m_axi_in_47_AWID,
  m_axi_in_47_AWLEN,
  m_axi_in_47_AWLOCK,
  m_axi_in_47_AWPROT,
  m_axi_in_47_AWQOS,
  m_axi_in_47_AWREADY,
  m_axi_in_47_AWSIZE,
  m_axi_in_47_AWVALID,
  m_axi_in_47_BID,
  m_axi_in_47_BREADY,
  m_axi_in_47_BRESP,
  m_axi_in_47_BVALID,
  m_axi_in_47_RDATA,
  m_axi_in_47_RID,
  m_axi_in_47_RLAST,
  m_axi_in_47_RREADY,
  m_axi_in_47_RRESP,
  m_axi_in_47_RVALID,
  m_axi_in_47_WDATA,
  m_axi_in_47_WLAST,
  m_axi_in_47_WREADY,
  m_axi_in_47_WSTRB,
  m_axi_in_47_WVALID,
  m_axi_in_48_ARADDR,
  m_axi_in_48_ARBURST,
  m_axi_in_48_ARCACHE,
  m_axi_in_48_ARID,
  m_axi_in_48_ARLEN,
  m_axi_in_48_ARLOCK,
  m_axi_in_48_ARPROT,
  m_axi_in_48_ARQOS,
  m_axi_in_48_ARREADY,
  m_axi_in_48_ARSIZE,
  m_axi_in_48_ARVALID,
  m_axi_in_48_AWADDR,
  m_axi_in_48_AWBURST,
  m_axi_in_48_AWCACHE,
  m_axi_in_48_AWID,
  m_axi_in_48_AWLEN,
  m_axi_in_48_AWLOCK,
  m_axi_in_48_AWPROT,
  m_axi_in_48_AWQOS,
  m_axi_in_48_AWREADY,
  m_axi_in_48_AWSIZE,
  m_axi_in_48_AWVALID,
  m_axi_in_48_BID,
  m_axi_in_48_BREADY,
  m_axi_in_48_BRESP,
  m_axi_in_48_BVALID,
  m_axi_in_48_RDATA,
  m_axi_in_48_RID,
  m_axi_in_48_RLAST,
  m_axi_in_48_RREADY,
  m_axi_in_48_RRESP,
  m_axi_in_48_RVALID,
  m_axi_in_48_WDATA,
  m_axi_in_48_WLAST,
  m_axi_in_48_WREADY,
  m_axi_in_48_WSTRB,
  m_axi_in_48_WVALID,
  m_axi_in_49_ARADDR,
  m_axi_in_49_ARBURST,
  m_axi_in_49_ARCACHE,
  m_axi_in_49_ARID,
  m_axi_in_49_ARLEN,
  m_axi_in_49_ARLOCK,
  m_axi_in_49_ARPROT,
  m_axi_in_49_ARQOS,
  m_axi_in_49_ARREADY,
  m_axi_in_49_ARSIZE,
  m_axi_in_49_ARVALID,
  m_axi_in_49_AWADDR,
  m_axi_in_49_AWBURST,
  m_axi_in_49_AWCACHE,
  m_axi_in_49_AWID,
  m_axi_in_49_AWLEN,
  m_axi_in_49_AWLOCK,
  m_axi_in_49_AWPROT,
  m_axi_in_49_AWQOS,
  m_axi_in_49_AWREADY,
  m_axi_in_49_AWSIZE,
  m_axi_in_49_AWVALID,
  m_axi_in_49_BID,
  m_axi_in_49_BREADY,
  m_axi_in_49_BRESP,
  m_axi_in_49_BVALID,
  m_axi_in_49_RDATA,
  m_axi_in_49_RID,
  m_axi_in_49_RLAST,
  m_axi_in_49_RREADY,
  m_axi_in_49_RRESP,
  m_axi_in_49_RVALID,
  m_axi_in_49_WDATA,
  m_axi_in_49_WLAST,
  m_axi_in_49_WREADY,
  m_axi_in_49_WSTRB,
  m_axi_in_49_WVALID,
  m_axi_in_5_ARADDR,
  m_axi_in_5_ARBURST,
  m_axi_in_5_ARCACHE,
  m_axi_in_5_ARID,
  m_axi_in_5_ARLEN,
  m_axi_in_5_ARLOCK,
  m_axi_in_5_ARPROT,
  m_axi_in_5_ARQOS,
  m_axi_in_5_ARREADY,
  m_axi_in_5_ARSIZE,
  m_axi_in_5_ARVALID,
  m_axi_in_5_AWADDR,
  m_axi_in_5_AWBURST,
  m_axi_in_5_AWCACHE,
  m_axi_in_5_AWID,
  m_axi_in_5_AWLEN,
  m_axi_in_5_AWLOCK,
  m_axi_in_5_AWPROT,
  m_axi_in_5_AWQOS,
  m_axi_in_5_AWREADY,
  m_axi_in_5_AWSIZE,
  m_axi_in_5_AWVALID,
  m_axi_in_5_BID,
  m_axi_in_5_BREADY,
  m_axi_in_5_BRESP,
  m_axi_in_5_BVALID,
  m_axi_in_5_RDATA,
  m_axi_in_5_RID,
  m_axi_in_5_RLAST,
  m_axi_in_5_RREADY,
  m_axi_in_5_RRESP,
  m_axi_in_5_RVALID,
  m_axi_in_5_WDATA,
  m_axi_in_5_WLAST,
  m_axi_in_5_WREADY,
  m_axi_in_5_WSTRB,
  m_axi_in_5_WVALID,
  m_axi_in_50_ARADDR,
  m_axi_in_50_ARBURST,
  m_axi_in_50_ARCACHE,
  m_axi_in_50_ARID,
  m_axi_in_50_ARLEN,
  m_axi_in_50_ARLOCK,
  m_axi_in_50_ARPROT,
  m_axi_in_50_ARQOS,
  m_axi_in_50_ARREADY,
  m_axi_in_50_ARSIZE,
  m_axi_in_50_ARVALID,
  m_axi_in_50_AWADDR,
  m_axi_in_50_AWBURST,
  m_axi_in_50_AWCACHE,
  m_axi_in_50_AWID,
  m_axi_in_50_AWLEN,
  m_axi_in_50_AWLOCK,
  m_axi_in_50_AWPROT,
  m_axi_in_50_AWQOS,
  m_axi_in_50_AWREADY,
  m_axi_in_50_AWSIZE,
  m_axi_in_50_AWVALID,
  m_axi_in_50_BID,
  m_axi_in_50_BREADY,
  m_axi_in_50_BRESP,
  m_axi_in_50_BVALID,
  m_axi_in_50_RDATA,
  m_axi_in_50_RID,
  m_axi_in_50_RLAST,
  m_axi_in_50_RREADY,
  m_axi_in_50_RRESP,
  m_axi_in_50_RVALID,
  m_axi_in_50_WDATA,
  m_axi_in_50_WLAST,
  m_axi_in_50_WREADY,
  m_axi_in_50_WSTRB,
  m_axi_in_50_WVALID,
  m_axi_in_51_ARADDR,
  m_axi_in_51_ARBURST,
  m_axi_in_51_ARCACHE,
  m_axi_in_51_ARID,
  m_axi_in_51_ARLEN,
  m_axi_in_51_ARLOCK,
  m_axi_in_51_ARPROT,
  m_axi_in_51_ARQOS,
  m_axi_in_51_ARREADY,
  m_axi_in_51_ARSIZE,
  m_axi_in_51_ARVALID,
  m_axi_in_51_AWADDR,
  m_axi_in_51_AWBURST,
  m_axi_in_51_AWCACHE,
  m_axi_in_51_AWID,
  m_axi_in_51_AWLEN,
  m_axi_in_51_AWLOCK,
  m_axi_in_51_AWPROT,
  m_axi_in_51_AWQOS,
  m_axi_in_51_AWREADY,
  m_axi_in_51_AWSIZE,
  m_axi_in_51_AWVALID,
  m_axi_in_51_BID,
  m_axi_in_51_BREADY,
  m_axi_in_51_BRESP,
  m_axi_in_51_BVALID,
  m_axi_in_51_RDATA,
  m_axi_in_51_RID,
  m_axi_in_51_RLAST,
  m_axi_in_51_RREADY,
  m_axi_in_51_RRESP,
  m_axi_in_51_RVALID,
  m_axi_in_51_WDATA,
  m_axi_in_51_WLAST,
  m_axi_in_51_WREADY,
  m_axi_in_51_WSTRB,
  m_axi_in_51_WVALID,
  m_axi_in_52_ARADDR,
  m_axi_in_52_ARBURST,
  m_axi_in_52_ARCACHE,
  m_axi_in_52_ARID,
  m_axi_in_52_ARLEN,
  m_axi_in_52_ARLOCK,
  m_axi_in_52_ARPROT,
  m_axi_in_52_ARQOS,
  m_axi_in_52_ARREADY,
  m_axi_in_52_ARSIZE,
  m_axi_in_52_ARVALID,
  m_axi_in_52_AWADDR,
  m_axi_in_52_AWBURST,
  m_axi_in_52_AWCACHE,
  m_axi_in_52_AWID,
  m_axi_in_52_AWLEN,
  m_axi_in_52_AWLOCK,
  m_axi_in_52_AWPROT,
  m_axi_in_52_AWQOS,
  m_axi_in_52_AWREADY,
  m_axi_in_52_AWSIZE,
  m_axi_in_52_AWVALID,
  m_axi_in_52_BID,
  m_axi_in_52_BREADY,
  m_axi_in_52_BRESP,
  m_axi_in_52_BVALID,
  m_axi_in_52_RDATA,
  m_axi_in_52_RID,
  m_axi_in_52_RLAST,
  m_axi_in_52_RREADY,
  m_axi_in_52_RRESP,
  m_axi_in_52_RVALID,
  m_axi_in_52_WDATA,
  m_axi_in_52_WLAST,
  m_axi_in_52_WREADY,
  m_axi_in_52_WSTRB,
  m_axi_in_52_WVALID,
  m_axi_in_53_ARADDR,
  m_axi_in_53_ARBURST,
  m_axi_in_53_ARCACHE,
  m_axi_in_53_ARID,
  m_axi_in_53_ARLEN,
  m_axi_in_53_ARLOCK,
  m_axi_in_53_ARPROT,
  m_axi_in_53_ARQOS,
  m_axi_in_53_ARREADY,
  m_axi_in_53_ARSIZE,
  m_axi_in_53_ARVALID,
  m_axi_in_53_AWADDR,
  m_axi_in_53_AWBURST,
  m_axi_in_53_AWCACHE,
  m_axi_in_53_AWID,
  m_axi_in_53_AWLEN,
  m_axi_in_53_AWLOCK,
  m_axi_in_53_AWPROT,
  m_axi_in_53_AWQOS,
  m_axi_in_53_AWREADY,
  m_axi_in_53_AWSIZE,
  m_axi_in_53_AWVALID,
  m_axi_in_53_BID,
  m_axi_in_53_BREADY,
  m_axi_in_53_BRESP,
  m_axi_in_53_BVALID,
  m_axi_in_53_RDATA,
  m_axi_in_53_RID,
  m_axi_in_53_RLAST,
  m_axi_in_53_RREADY,
  m_axi_in_53_RRESP,
  m_axi_in_53_RVALID,
  m_axi_in_53_WDATA,
  m_axi_in_53_WLAST,
  m_axi_in_53_WREADY,
  m_axi_in_53_WSTRB,
  m_axi_in_53_WVALID,
  m_axi_in_6_ARADDR,
  m_axi_in_6_ARBURST,
  m_axi_in_6_ARCACHE,
  m_axi_in_6_ARID,
  m_axi_in_6_ARLEN,
  m_axi_in_6_ARLOCK,
  m_axi_in_6_ARPROT,
  m_axi_in_6_ARQOS,
  m_axi_in_6_ARREADY,
  m_axi_in_6_ARSIZE,
  m_axi_in_6_ARVALID,
  m_axi_in_6_AWADDR,
  m_axi_in_6_AWBURST,
  m_axi_in_6_AWCACHE,
  m_axi_in_6_AWID,
  m_axi_in_6_AWLEN,
  m_axi_in_6_AWLOCK,
  m_axi_in_6_AWPROT,
  m_axi_in_6_AWQOS,
  m_axi_in_6_AWREADY,
  m_axi_in_6_AWSIZE,
  m_axi_in_6_AWVALID,
  m_axi_in_6_BID,
  m_axi_in_6_BREADY,
  m_axi_in_6_BRESP,
  m_axi_in_6_BVALID,
  m_axi_in_6_RDATA,
  m_axi_in_6_RID,
  m_axi_in_6_RLAST,
  m_axi_in_6_RREADY,
  m_axi_in_6_RRESP,
  m_axi_in_6_RVALID,
  m_axi_in_6_WDATA,
  m_axi_in_6_WLAST,
  m_axi_in_6_WREADY,
  m_axi_in_6_WSTRB,
  m_axi_in_6_WVALID,
  m_axi_in_7_ARADDR,
  m_axi_in_7_ARBURST,
  m_axi_in_7_ARCACHE,
  m_axi_in_7_ARID,
  m_axi_in_7_ARLEN,
  m_axi_in_7_ARLOCK,
  m_axi_in_7_ARPROT,
  m_axi_in_7_ARQOS,
  m_axi_in_7_ARREADY,
  m_axi_in_7_ARSIZE,
  m_axi_in_7_ARVALID,
  m_axi_in_7_AWADDR,
  m_axi_in_7_AWBURST,
  m_axi_in_7_AWCACHE,
  m_axi_in_7_AWID,
  m_axi_in_7_AWLEN,
  m_axi_in_7_AWLOCK,
  m_axi_in_7_AWPROT,
  m_axi_in_7_AWQOS,
  m_axi_in_7_AWREADY,
  m_axi_in_7_AWSIZE,
  m_axi_in_7_AWVALID,
  m_axi_in_7_BID,
  m_axi_in_7_BREADY,
  m_axi_in_7_BRESP,
  m_axi_in_7_BVALID,
  m_axi_in_7_RDATA,
  m_axi_in_7_RID,
  m_axi_in_7_RLAST,
  m_axi_in_7_RREADY,
  m_axi_in_7_RRESP,
  m_axi_in_7_RVALID,
  m_axi_in_7_WDATA,
  m_axi_in_7_WLAST,
  m_axi_in_7_WREADY,
  m_axi_in_7_WSTRB,
  m_axi_in_7_WVALID,
  m_axi_in_8_ARADDR,
  m_axi_in_8_ARBURST,
  m_axi_in_8_ARCACHE,
  m_axi_in_8_ARID,
  m_axi_in_8_ARLEN,
  m_axi_in_8_ARLOCK,
  m_axi_in_8_ARPROT,
  m_axi_in_8_ARQOS,
  m_axi_in_8_ARREADY,
  m_axi_in_8_ARSIZE,
  m_axi_in_8_ARVALID,
  m_axi_in_8_AWADDR,
  m_axi_in_8_AWBURST,
  m_axi_in_8_AWCACHE,
  m_axi_in_8_AWID,
  m_axi_in_8_AWLEN,
  m_axi_in_8_AWLOCK,
  m_axi_in_8_AWPROT,
  m_axi_in_8_AWQOS,
  m_axi_in_8_AWREADY,
  m_axi_in_8_AWSIZE,
  m_axi_in_8_AWVALID,
  m_axi_in_8_BID,
  m_axi_in_8_BREADY,
  m_axi_in_8_BRESP,
  m_axi_in_8_BVALID,
  m_axi_in_8_RDATA,
  m_axi_in_8_RID,
  m_axi_in_8_RLAST,
  m_axi_in_8_RREADY,
  m_axi_in_8_RRESP,
  m_axi_in_8_RVALID,
  m_axi_in_8_WDATA,
  m_axi_in_8_WLAST,
  m_axi_in_8_WREADY,
  m_axi_in_8_WSTRB,
  m_axi_in_8_WVALID,
  m_axi_in_9_ARADDR,
  m_axi_in_9_ARBURST,
  m_axi_in_9_ARCACHE,
  m_axi_in_9_ARID,
  m_axi_in_9_ARLEN,
  m_axi_in_9_ARLOCK,
  m_axi_in_9_ARPROT,
  m_axi_in_9_ARQOS,
  m_axi_in_9_ARREADY,
  m_axi_in_9_ARSIZE,
  m_axi_in_9_ARVALID,
  m_axi_in_9_AWADDR,
  m_axi_in_9_AWBURST,
  m_axi_in_9_AWCACHE,
  m_axi_in_9_AWID,
  m_axi_in_9_AWLEN,
  m_axi_in_9_AWLOCK,
  m_axi_in_9_AWPROT,
  m_axi_in_9_AWQOS,
  m_axi_in_9_AWREADY,
  m_axi_in_9_AWSIZE,
  m_axi_in_9_AWVALID,
  m_axi_in_9_BID,
  m_axi_in_9_BREADY,
  m_axi_in_9_BRESP,
  m_axi_in_9_BVALID,
  m_axi_in_9_RDATA,
  m_axi_in_9_RID,
  m_axi_in_9_RLAST,
  m_axi_in_9_RREADY,
  m_axi_in_9_RRESP,
  m_axi_in_9_RVALID,
  m_axi_in_9_WDATA,
  m_axi_in_9_WLAST,
  m_axi_in_9_WREADY,
  m_axi_in_9_WSTRB,
  m_axi_in_9_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 10;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [63:0] m_axi_L4_out_dist_ARADDR;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [1:0] m_axi_L4_out_dist_ARBURST;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [3:0] m_axi_L4_out_dist_ARCACHE;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [0:0] m_axi_L4_out_dist_ARID;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [7:0] m_axi_L4_out_dist_ARLEN;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output m_axi_L4_out_dist_ARLOCK;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [2:0] m_axi_L4_out_dist_ARPROT;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [3:0] m_axi_L4_out_dist_ARQOS;
  (* RS_HS = "m_axi_L4_out_dist_AR.ready" *)input m_axi_L4_out_dist_ARREADY;
  (* RS_HS = "m_axi_L4_out_dist_AR.data" *)output [2:0] m_axi_L4_out_dist_ARSIZE;
  (* RS_HS = "m_axi_L4_out_dist_AR.valid" *)output m_axi_L4_out_dist_ARVALID;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [63:0] m_axi_L4_out_dist_AWADDR;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [1:0] m_axi_L4_out_dist_AWBURST;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [3:0] m_axi_L4_out_dist_AWCACHE;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [0:0] m_axi_L4_out_dist_AWID;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [7:0] m_axi_L4_out_dist_AWLEN;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output m_axi_L4_out_dist_AWLOCK;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [2:0] m_axi_L4_out_dist_AWPROT;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [3:0] m_axi_L4_out_dist_AWQOS;
  (* RS_HS = "m_axi_L4_out_dist_AW.ready" *)input m_axi_L4_out_dist_AWREADY;
  (* RS_HS = "m_axi_L4_out_dist_AW.data" *)output [2:0] m_axi_L4_out_dist_AWSIZE;
  (* RS_HS = "m_axi_L4_out_dist_AW.valid" *)output m_axi_L4_out_dist_AWVALID;
  (* RS_HS = "m_axi_L4_out_dist_B.data" *)input [0:0] m_axi_L4_out_dist_BID;
  (* RS_HS = "m_axi_L4_out_dist_B.ready" *)output m_axi_L4_out_dist_BREADY;
  (* RS_HS = "m_axi_L4_out_dist_B.data" *)input [1:0] m_axi_L4_out_dist_BRESP;
  (* RS_HS = "m_axi_L4_out_dist_B.valid" *)input m_axi_L4_out_dist_BVALID;
  (* RS_HS = "m_axi_L4_out_dist_R.data" *)input [31:0] m_axi_L4_out_dist_RDATA;
  (* RS_HS = "m_axi_L4_out_dist_R.data" *)input [0:0] m_axi_L4_out_dist_RID;
  (* RS_HS = "m_axi_L4_out_dist_R.data" *)input m_axi_L4_out_dist_RLAST;
  (* RS_HS = "m_axi_L4_out_dist_R.ready" *)output m_axi_L4_out_dist_RREADY;
  (* RS_HS = "m_axi_L4_out_dist_R.data" *)input [1:0] m_axi_L4_out_dist_RRESP;
  (* RS_HS = "m_axi_L4_out_dist_R.valid" *)input m_axi_L4_out_dist_RVALID;
  (* RS_HS = "m_axi_L4_out_dist_W.data" *)output [31:0] m_axi_L4_out_dist_WDATA;
  (* RS_HS = "m_axi_L4_out_dist_W.data" *)output m_axi_L4_out_dist_WLAST;
  (* RS_HS = "m_axi_L4_out_dist_W.ready" *)input m_axi_L4_out_dist_WREADY;
  (* RS_HS = "m_axi_L4_out_dist_W.data" *)output [3:0] m_axi_L4_out_dist_WSTRB;
  (* RS_HS = "m_axi_L4_out_dist_W.valid" *)output m_axi_L4_out_dist_WVALID;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [63:0] m_axi_L4_out_id_ARADDR;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [1:0] m_axi_L4_out_id_ARBURST;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [3:0] m_axi_L4_out_id_ARCACHE;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [0:0] m_axi_L4_out_id_ARID;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [7:0] m_axi_L4_out_id_ARLEN;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output m_axi_L4_out_id_ARLOCK;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [2:0] m_axi_L4_out_id_ARPROT;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [3:0] m_axi_L4_out_id_ARQOS;
  (* RS_HS = "m_axi_L4_out_id_AR.ready" *)input m_axi_L4_out_id_ARREADY;
  (* RS_HS = "m_axi_L4_out_id_AR.data" *)output [2:0] m_axi_L4_out_id_ARSIZE;
  (* RS_HS = "m_axi_L4_out_id_AR.valid" *)output m_axi_L4_out_id_ARVALID;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [63:0] m_axi_L4_out_id_AWADDR;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [1:0] m_axi_L4_out_id_AWBURST;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [3:0] m_axi_L4_out_id_AWCACHE;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [0:0] m_axi_L4_out_id_AWID;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [7:0] m_axi_L4_out_id_AWLEN;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output m_axi_L4_out_id_AWLOCK;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [2:0] m_axi_L4_out_id_AWPROT;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [3:0] m_axi_L4_out_id_AWQOS;
  (* RS_HS = "m_axi_L4_out_id_AW.ready" *)input m_axi_L4_out_id_AWREADY;
  (* RS_HS = "m_axi_L4_out_id_AW.data" *)output [2:0] m_axi_L4_out_id_AWSIZE;
  (* RS_HS = "m_axi_L4_out_id_AW.valid" *)output m_axi_L4_out_id_AWVALID;
  (* RS_HS = "m_axi_L4_out_id_B.data" *)input [0:0] m_axi_L4_out_id_BID;
  (* RS_HS = "m_axi_L4_out_id_B.ready" *)output m_axi_L4_out_id_BREADY;
  (* RS_HS = "m_axi_L4_out_id_B.data" *)input [1:0] m_axi_L4_out_id_BRESP;
  (* RS_HS = "m_axi_L4_out_id_B.valid" *)input m_axi_L4_out_id_BVALID;
  (* RS_HS = "m_axi_L4_out_id_R.data" *)input [31:0] m_axi_L4_out_id_RDATA;
  (* RS_HS = "m_axi_L4_out_id_R.data" *)input [0:0] m_axi_L4_out_id_RID;
  (* RS_HS = "m_axi_L4_out_id_R.data" *)input m_axi_L4_out_id_RLAST;
  (* RS_HS = "m_axi_L4_out_id_R.ready" *)output m_axi_L4_out_id_RREADY;
  (* RS_HS = "m_axi_L4_out_id_R.data" *)input [1:0] m_axi_L4_out_id_RRESP;
  (* RS_HS = "m_axi_L4_out_id_R.valid" *)input m_axi_L4_out_id_RVALID;
  (* RS_HS = "m_axi_L4_out_id_W.data" *)output [31:0] m_axi_L4_out_id_WDATA;
  (* RS_HS = "m_axi_L4_out_id_W.data" *)output m_axi_L4_out_id_WLAST;
  (* RS_HS = "m_axi_L4_out_id_W.ready" *)input m_axi_L4_out_id_WREADY;
  (* RS_HS = "m_axi_L4_out_id_W.data" *)output [3:0] m_axi_L4_out_id_WSTRB;
  (* RS_HS = "m_axi_L4_out_id_W.valid" *)output m_axi_L4_out_id_WVALID;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [63:0] m_axi_in_0_ARADDR;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [1:0] m_axi_in_0_ARBURST;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [3:0] m_axi_in_0_ARCACHE;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [0:0] m_axi_in_0_ARID;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [7:0] m_axi_in_0_ARLEN;
  (* RS_HS = "m_axi_in_0_AR.data" *)output m_axi_in_0_ARLOCK;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [2:0] m_axi_in_0_ARPROT;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [3:0] m_axi_in_0_ARQOS;
  (* RS_HS = "m_axi_in_0_AR.ready" *)input m_axi_in_0_ARREADY;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [2:0] m_axi_in_0_ARSIZE;
  (* RS_HS = "m_axi_in_0_AR.valid" *)output m_axi_in_0_ARVALID;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [63:0] m_axi_in_0_AWADDR;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [1:0] m_axi_in_0_AWBURST;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [3:0] m_axi_in_0_AWCACHE;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [0:0] m_axi_in_0_AWID;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [7:0] m_axi_in_0_AWLEN;
  (* RS_HS = "m_axi_in_0_AW.data" *)output m_axi_in_0_AWLOCK;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [2:0] m_axi_in_0_AWPROT;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [3:0] m_axi_in_0_AWQOS;
  (* RS_HS = "m_axi_in_0_AW.ready" *)input m_axi_in_0_AWREADY;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [2:0] m_axi_in_0_AWSIZE;
  (* RS_HS = "m_axi_in_0_AW.valid" *)output m_axi_in_0_AWVALID;
  (* RS_HS = "m_axi_in_0_B.data" *)input [0:0] m_axi_in_0_BID;
  (* RS_HS = "m_axi_in_0_B.ready" *)output m_axi_in_0_BREADY;
  (* RS_HS = "m_axi_in_0_B.data" *)input [1:0] m_axi_in_0_BRESP;
  (* RS_HS = "m_axi_in_0_B.valid" *)input m_axi_in_0_BVALID;
  (* RS_HS = "m_axi_in_0_R.data" *)input [255:0] m_axi_in_0_RDATA;
  (* RS_HS = "m_axi_in_0_R.data" *)input [0:0] m_axi_in_0_RID;
  (* RS_HS = "m_axi_in_0_R.data" *)input m_axi_in_0_RLAST;
  (* RS_HS = "m_axi_in_0_R.ready" *)output m_axi_in_0_RREADY;
  (* RS_HS = "m_axi_in_0_R.data" *)input [1:0] m_axi_in_0_RRESP;
  (* RS_HS = "m_axi_in_0_R.valid" *)input m_axi_in_0_RVALID;
  (* RS_HS = "m_axi_in_0_W.data" *)output [255:0] m_axi_in_0_WDATA;
  (* RS_HS = "m_axi_in_0_W.data" *)output m_axi_in_0_WLAST;
  (* RS_HS = "m_axi_in_0_W.ready" *)input m_axi_in_0_WREADY;
  (* RS_HS = "m_axi_in_0_W.data" *)output [31:0] m_axi_in_0_WSTRB;
  (* RS_HS = "m_axi_in_0_W.valid" *)output m_axi_in_0_WVALID;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [63:0] m_axi_in_1_ARADDR;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [1:0] m_axi_in_1_ARBURST;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [3:0] m_axi_in_1_ARCACHE;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [0:0] m_axi_in_1_ARID;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [7:0] m_axi_in_1_ARLEN;
  (* RS_HS = "m_axi_in_1_AR.data" *)output m_axi_in_1_ARLOCK;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [2:0] m_axi_in_1_ARPROT;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [3:0] m_axi_in_1_ARQOS;
  (* RS_HS = "m_axi_in_1_AR.ready" *)input m_axi_in_1_ARREADY;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [2:0] m_axi_in_1_ARSIZE;
  (* RS_HS = "m_axi_in_1_AR.valid" *)output m_axi_in_1_ARVALID;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [63:0] m_axi_in_1_AWADDR;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [1:0] m_axi_in_1_AWBURST;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [3:0] m_axi_in_1_AWCACHE;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [0:0] m_axi_in_1_AWID;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [7:0] m_axi_in_1_AWLEN;
  (* RS_HS = "m_axi_in_1_AW.data" *)output m_axi_in_1_AWLOCK;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [2:0] m_axi_in_1_AWPROT;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [3:0] m_axi_in_1_AWQOS;
  (* RS_HS = "m_axi_in_1_AW.ready" *)input m_axi_in_1_AWREADY;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [2:0] m_axi_in_1_AWSIZE;
  (* RS_HS = "m_axi_in_1_AW.valid" *)output m_axi_in_1_AWVALID;
  (* RS_HS = "m_axi_in_1_B.data" *)input [0:0] m_axi_in_1_BID;
  (* RS_HS = "m_axi_in_1_B.ready" *)output m_axi_in_1_BREADY;
  (* RS_HS = "m_axi_in_1_B.data" *)input [1:0] m_axi_in_1_BRESP;
  (* RS_HS = "m_axi_in_1_B.valid" *)input m_axi_in_1_BVALID;
  (* RS_HS = "m_axi_in_1_R.data" *)input [255:0] m_axi_in_1_RDATA;
  (* RS_HS = "m_axi_in_1_R.data" *)input [0:0] m_axi_in_1_RID;
  (* RS_HS = "m_axi_in_1_R.data" *)input m_axi_in_1_RLAST;
  (* RS_HS = "m_axi_in_1_R.ready" *)output m_axi_in_1_RREADY;
  (* RS_HS = "m_axi_in_1_R.data" *)input [1:0] m_axi_in_1_RRESP;
  (* RS_HS = "m_axi_in_1_R.valid" *)input m_axi_in_1_RVALID;
  (* RS_HS = "m_axi_in_1_W.data" *)output [255:0] m_axi_in_1_WDATA;
  (* RS_HS = "m_axi_in_1_W.data" *)output m_axi_in_1_WLAST;
  (* RS_HS = "m_axi_in_1_W.ready" *)input m_axi_in_1_WREADY;
  (* RS_HS = "m_axi_in_1_W.data" *)output [31:0] m_axi_in_1_WSTRB;
  (* RS_HS = "m_axi_in_1_W.valid" *)output m_axi_in_1_WVALID;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [63:0] m_axi_in_10_ARADDR;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [1:0] m_axi_in_10_ARBURST;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [3:0] m_axi_in_10_ARCACHE;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [0:0] m_axi_in_10_ARID;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [7:0] m_axi_in_10_ARLEN;
  (* RS_HS = "m_axi_in_10_AR.data" *)output m_axi_in_10_ARLOCK;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [2:0] m_axi_in_10_ARPROT;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [3:0] m_axi_in_10_ARQOS;
  (* RS_HS = "m_axi_in_10_AR.ready" *)input m_axi_in_10_ARREADY;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [2:0] m_axi_in_10_ARSIZE;
  (* RS_HS = "m_axi_in_10_AR.valid" *)output m_axi_in_10_ARVALID;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [63:0] m_axi_in_10_AWADDR;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [1:0] m_axi_in_10_AWBURST;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [3:0] m_axi_in_10_AWCACHE;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [0:0] m_axi_in_10_AWID;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [7:0] m_axi_in_10_AWLEN;
  (* RS_HS = "m_axi_in_10_AW.data" *)output m_axi_in_10_AWLOCK;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [2:0] m_axi_in_10_AWPROT;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [3:0] m_axi_in_10_AWQOS;
  (* RS_HS = "m_axi_in_10_AW.ready" *)input m_axi_in_10_AWREADY;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [2:0] m_axi_in_10_AWSIZE;
  (* RS_HS = "m_axi_in_10_AW.valid" *)output m_axi_in_10_AWVALID;
  (* RS_HS = "m_axi_in_10_B.data" *)input [0:0] m_axi_in_10_BID;
  (* RS_HS = "m_axi_in_10_B.ready" *)output m_axi_in_10_BREADY;
  (* RS_HS = "m_axi_in_10_B.data" *)input [1:0] m_axi_in_10_BRESP;
  (* RS_HS = "m_axi_in_10_B.valid" *)input m_axi_in_10_BVALID;
  (* RS_HS = "m_axi_in_10_R.data" *)input [255:0] m_axi_in_10_RDATA;
  (* RS_HS = "m_axi_in_10_R.data" *)input [0:0] m_axi_in_10_RID;
  (* RS_HS = "m_axi_in_10_R.data" *)input m_axi_in_10_RLAST;
  (* RS_HS = "m_axi_in_10_R.ready" *)output m_axi_in_10_RREADY;
  (* RS_HS = "m_axi_in_10_R.data" *)input [1:0] m_axi_in_10_RRESP;
  (* RS_HS = "m_axi_in_10_R.valid" *)input m_axi_in_10_RVALID;
  (* RS_HS = "m_axi_in_10_W.data" *)output [255:0] m_axi_in_10_WDATA;
  (* RS_HS = "m_axi_in_10_W.data" *)output m_axi_in_10_WLAST;
  (* RS_HS = "m_axi_in_10_W.ready" *)input m_axi_in_10_WREADY;
  (* RS_HS = "m_axi_in_10_W.data" *)output [31:0] m_axi_in_10_WSTRB;
  (* RS_HS = "m_axi_in_10_W.valid" *)output m_axi_in_10_WVALID;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [63:0] m_axi_in_11_ARADDR;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [1:0] m_axi_in_11_ARBURST;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [3:0] m_axi_in_11_ARCACHE;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [0:0] m_axi_in_11_ARID;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [7:0] m_axi_in_11_ARLEN;
  (* RS_HS = "m_axi_in_11_AR.data" *)output m_axi_in_11_ARLOCK;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [2:0] m_axi_in_11_ARPROT;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [3:0] m_axi_in_11_ARQOS;
  (* RS_HS = "m_axi_in_11_AR.ready" *)input m_axi_in_11_ARREADY;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [2:0] m_axi_in_11_ARSIZE;
  (* RS_HS = "m_axi_in_11_AR.valid" *)output m_axi_in_11_ARVALID;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [63:0] m_axi_in_11_AWADDR;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [1:0] m_axi_in_11_AWBURST;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [3:0] m_axi_in_11_AWCACHE;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [0:0] m_axi_in_11_AWID;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [7:0] m_axi_in_11_AWLEN;
  (* RS_HS = "m_axi_in_11_AW.data" *)output m_axi_in_11_AWLOCK;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [2:0] m_axi_in_11_AWPROT;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [3:0] m_axi_in_11_AWQOS;
  (* RS_HS = "m_axi_in_11_AW.ready" *)input m_axi_in_11_AWREADY;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [2:0] m_axi_in_11_AWSIZE;
  (* RS_HS = "m_axi_in_11_AW.valid" *)output m_axi_in_11_AWVALID;
  (* RS_HS = "m_axi_in_11_B.data" *)input [0:0] m_axi_in_11_BID;
  (* RS_HS = "m_axi_in_11_B.ready" *)output m_axi_in_11_BREADY;
  (* RS_HS = "m_axi_in_11_B.data" *)input [1:0] m_axi_in_11_BRESP;
  (* RS_HS = "m_axi_in_11_B.valid" *)input m_axi_in_11_BVALID;
  (* RS_HS = "m_axi_in_11_R.data" *)input [255:0] m_axi_in_11_RDATA;
  (* RS_HS = "m_axi_in_11_R.data" *)input [0:0] m_axi_in_11_RID;
  (* RS_HS = "m_axi_in_11_R.data" *)input m_axi_in_11_RLAST;
  (* RS_HS = "m_axi_in_11_R.ready" *)output m_axi_in_11_RREADY;
  (* RS_HS = "m_axi_in_11_R.data" *)input [1:0] m_axi_in_11_RRESP;
  (* RS_HS = "m_axi_in_11_R.valid" *)input m_axi_in_11_RVALID;
  (* RS_HS = "m_axi_in_11_W.data" *)output [255:0] m_axi_in_11_WDATA;
  (* RS_HS = "m_axi_in_11_W.data" *)output m_axi_in_11_WLAST;
  (* RS_HS = "m_axi_in_11_W.ready" *)input m_axi_in_11_WREADY;
  (* RS_HS = "m_axi_in_11_W.data" *)output [31:0] m_axi_in_11_WSTRB;
  (* RS_HS = "m_axi_in_11_W.valid" *)output m_axi_in_11_WVALID;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [63:0] m_axi_in_12_ARADDR;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [1:0] m_axi_in_12_ARBURST;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [3:0] m_axi_in_12_ARCACHE;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [0:0] m_axi_in_12_ARID;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [7:0] m_axi_in_12_ARLEN;
  (* RS_HS = "m_axi_in_12_AR.data" *)output m_axi_in_12_ARLOCK;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [2:0] m_axi_in_12_ARPROT;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [3:0] m_axi_in_12_ARQOS;
  (* RS_HS = "m_axi_in_12_AR.ready" *)input m_axi_in_12_ARREADY;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [2:0] m_axi_in_12_ARSIZE;
  (* RS_HS = "m_axi_in_12_AR.valid" *)output m_axi_in_12_ARVALID;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [63:0] m_axi_in_12_AWADDR;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [1:0] m_axi_in_12_AWBURST;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [3:0] m_axi_in_12_AWCACHE;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [0:0] m_axi_in_12_AWID;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [7:0] m_axi_in_12_AWLEN;
  (* RS_HS = "m_axi_in_12_AW.data" *)output m_axi_in_12_AWLOCK;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [2:0] m_axi_in_12_AWPROT;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [3:0] m_axi_in_12_AWQOS;
  (* RS_HS = "m_axi_in_12_AW.ready" *)input m_axi_in_12_AWREADY;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [2:0] m_axi_in_12_AWSIZE;
  (* RS_HS = "m_axi_in_12_AW.valid" *)output m_axi_in_12_AWVALID;
  (* RS_HS = "m_axi_in_12_B.data" *)input [0:0] m_axi_in_12_BID;
  (* RS_HS = "m_axi_in_12_B.ready" *)output m_axi_in_12_BREADY;
  (* RS_HS = "m_axi_in_12_B.data" *)input [1:0] m_axi_in_12_BRESP;
  (* RS_HS = "m_axi_in_12_B.valid" *)input m_axi_in_12_BVALID;
  (* RS_HS = "m_axi_in_12_R.data" *)input [255:0] m_axi_in_12_RDATA;
  (* RS_HS = "m_axi_in_12_R.data" *)input [0:0] m_axi_in_12_RID;
  (* RS_HS = "m_axi_in_12_R.data" *)input m_axi_in_12_RLAST;
  (* RS_HS = "m_axi_in_12_R.ready" *)output m_axi_in_12_RREADY;
  (* RS_HS = "m_axi_in_12_R.data" *)input [1:0] m_axi_in_12_RRESP;
  (* RS_HS = "m_axi_in_12_R.valid" *)input m_axi_in_12_RVALID;
  (* RS_HS = "m_axi_in_12_W.data" *)output [255:0] m_axi_in_12_WDATA;
  (* RS_HS = "m_axi_in_12_W.data" *)output m_axi_in_12_WLAST;
  (* RS_HS = "m_axi_in_12_W.ready" *)input m_axi_in_12_WREADY;
  (* RS_HS = "m_axi_in_12_W.data" *)output [31:0] m_axi_in_12_WSTRB;
  (* RS_HS = "m_axi_in_12_W.valid" *)output m_axi_in_12_WVALID;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [63:0] m_axi_in_13_ARADDR;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [1:0] m_axi_in_13_ARBURST;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [3:0] m_axi_in_13_ARCACHE;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [0:0] m_axi_in_13_ARID;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [7:0] m_axi_in_13_ARLEN;
  (* RS_HS = "m_axi_in_13_AR.data" *)output m_axi_in_13_ARLOCK;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [2:0] m_axi_in_13_ARPROT;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [3:0] m_axi_in_13_ARQOS;
  (* RS_HS = "m_axi_in_13_AR.ready" *)input m_axi_in_13_ARREADY;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [2:0] m_axi_in_13_ARSIZE;
  (* RS_HS = "m_axi_in_13_AR.valid" *)output m_axi_in_13_ARVALID;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [63:0] m_axi_in_13_AWADDR;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [1:0] m_axi_in_13_AWBURST;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [3:0] m_axi_in_13_AWCACHE;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [0:0] m_axi_in_13_AWID;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [7:0] m_axi_in_13_AWLEN;
  (* RS_HS = "m_axi_in_13_AW.data" *)output m_axi_in_13_AWLOCK;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [2:0] m_axi_in_13_AWPROT;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [3:0] m_axi_in_13_AWQOS;
  (* RS_HS = "m_axi_in_13_AW.ready" *)input m_axi_in_13_AWREADY;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [2:0] m_axi_in_13_AWSIZE;
  (* RS_HS = "m_axi_in_13_AW.valid" *)output m_axi_in_13_AWVALID;
  (* RS_HS = "m_axi_in_13_B.data" *)input [0:0] m_axi_in_13_BID;
  (* RS_HS = "m_axi_in_13_B.ready" *)output m_axi_in_13_BREADY;
  (* RS_HS = "m_axi_in_13_B.data" *)input [1:0] m_axi_in_13_BRESP;
  (* RS_HS = "m_axi_in_13_B.valid" *)input m_axi_in_13_BVALID;
  (* RS_HS = "m_axi_in_13_R.data" *)input [255:0] m_axi_in_13_RDATA;
  (* RS_HS = "m_axi_in_13_R.data" *)input [0:0] m_axi_in_13_RID;
  (* RS_HS = "m_axi_in_13_R.data" *)input m_axi_in_13_RLAST;
  (* RS_HS = "m_axi_in_13_R.ready" *)output m_axi_in_13_RREADY;
  (* RS_HS = "m_axi_in_13_R.data" *)input [1:0] m_axi_in_13_RRESP;
  (* RS_HS = "m_axi_in_13_R.valid" *)input m_axi_in_13_RVALID;
  (* RS_HS = "m_axi_in_13_W.data" *)output [255:0] m_axi_in_13_WDATA;
  (* RS_HS = "m_axi_in_13_W.data" *)output m_axi_in_13_WLAST;
  (* RS_HS = "m_axi_in_13_W.ready" *)input m_axi_in_13_WREADY;
  (* RS_HS = "m_axi_in_13_W.data" *)output [31:0] m_axi_in_13_WSTRB;
  (* RS_HS = "m_axi_in_13_W.valid" *)output m_axi_in_13_WVALID;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [63:0] m_axi_in_14_ARADDR;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [1:0] m_axi_in_14_ARBURST;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [3:0] m_axi_in_14_ARCACHE;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [0:0] m_axi_in_14_ARID;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [7:0] m_axi_in_14_ARLEN;
  (* RS_HS = "m_axi_in_14_AR.data" *)output m_axi_in_14_ARLOCK;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [2:0] m_axi_in_14_ARPROT;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [3:0] m_axi_in_14_ARQOS;
  (* RS_HS = "m_axi_in_14_AR.ready" *)input m_axi_in_14_ARREADY;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [2:0] m_axi_in_14_ARSIZE;
  (* RS_HS = "m_axi_in_14_AR.valid" *)output m_axi_in_14_ARVALID;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [63:0] m_axi_in_14_AWADDR;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [1:0] m_axi_in_14_AWBURST;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [3:0] m_axi_in_14_AWCACHE;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [0:0] m_axi_in_14_AWID;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [7:0] m_axi_in_14_AWLEN;
  (* RS_HS = "m_axi_in_14_AW.data" *)output m_axi_in_14_AWLOCK;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [2:0] m_axi_in_14_AWPROT;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [3:0] m_axi_in_14_AWQOS;
  (* RS_HS = "m_axi_in_14_AW.ready" *)input m_axi_in_14_AWREADY;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [2:0] m_axi_in_14_AWSIZE;
  (* RS_HS = "m_axi_in_14_AW.valid" *)output m_axi_in_14_AWVALID;
  (* RS_HS = "m_axi_in_14_B.data" *)input [0:0] m_axi_in_14_BID;
  (* RS_HS = "m_axi_in_14_B.ready" *)output m_axi_in_14_BREADY;
  (* RS_HS = "m_axi_in_14_B.data" *)input [1:0] m_axi_in_14_BRESP;
  (* RS_HS = "m_axi_in_14_B.valid" *)input m_axi_in_14_BVALID;
  (* RS_HS = "m_axi_in_14_R.data" *)input [255:0] m_axi_in_14_RDATA;
  (* RS_HS = "m_axi_in_14_R.data" *)input [0:0] m_axi_in_14_RID;
  (* RS_HS = "m_axi_in_14_R.data" *)input m_axi_in_14_RLAST;
  (* RS_HS = "m_axi_in_14_R.ready" *)output m_axi_in_14_RREADY;
  (* RS_HS = "m_axi_in_14_R.data" *)input [1:0] m_axi_in_14_RRESP;
  (* RS_HS = "m_axi_in_14_R.valid" *)input m_axi_in_14_RVALID;
  (* RS_HS = "m_axi_in_14_W.data" *)output [255:0] m_axi_in_14_WDATA;
  (* RS_HS = "m_axi_in_14_W.data" *)output m_axi_in_14_WLAST;
  (* RS_HS = "m_axi_in_14_W.ready" *)input m_axi_in_14_WREADY;
  (* RS_HS = "m_axi_in_14_W.data" *)output [31:0] m_axi_in_14_WSTRB;
  (* RS_HS = "m_axi_in_14_W.valid" *)output m_axi_in_14_WVALID;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [63:0] m_axi_in_15_ARADDR;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [1:0] m_axi_in_15_ARBURST;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [3:0] m_axi_in_15_ARCACHE;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [0:0] m_axi_in_15_ARID;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [7:0] m_axi_in_15_ARLEN;
  (* RS_HS = "m_axi_in_15_AR.data" *)output m_axi_in_15_ARLOCK;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [2:0] m_axi_in_15_ARPROT;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [3:0] m_axi_in_15_ARQOS;
  (* RS_HS = "m_axi_in_15_AR.ready" *)input m_axi_in_15_ARREADY;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [2:0] m_axi_in_15_ARSIZE;
  (* RS_HS = "m_axi_in_15_AR.valid" *)output m_axi_in_15_ARVALID;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [63:0] m_axi_in_15_AWADDR;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [1:0] m_axi_in_15_AWBURST;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [3:0] m_axi_in_15_AWCACHE;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [0:0] m_axi_in_15_AWID;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [7:0] m_axi_in_15_AWLEN;
  (* RS_HS = "m_axi_in_15_AW.data" *)output m_axi_in_15_AWLOCK;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [2:0] m_axi_in_15_AWPROT;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [3:0] m_axi_in_15_AWQOS;
  (* RS_HS = "m_axi_in_15_AW.ready" *)input m_axi_in_15_AWREADY;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [2:0] m_axi_in_15_AWSIZE;
  (* RS_HS = "m_axi_in_15_AW.valid" *)output m_axi_in_15_AWVALID;
  (* RS_HS = "m_axi_in_15_B.data" *)input [0:0] m_axi_in_15_BID;
  (* RS_HS = "m_axi_in_15_B.ready" *)output m_axi_in_15_BREADY;
  (* RS_HS = "m_axi_in_15_B.data" *)input [1:0] m_axi_in_15_BRESP;
  (* RS_HS = "m_axi_in_15_B.valid" *)input m_axi_in_15_BVALID;
  (* RS_HS = "m_axi_in_15_R.data" *)input [255:0] m_axi_in_15_RDATA;
  (* RS_HS = "m_axi_in_15_R.data" *)input [0:0] m_axi_in_15_RID;
  (* RS_HS = "m_axi_in_15_R.data" *)input m_axi_in_15_RLAST;
  (* RS_HS = "m_axi_in_15_R.ready" *)output m_axi_in_15_RREADY;
  (* RS_HS = "m_axi_in_15_R.data" *)input [1:0] m_axi_in_15_RRESP;
  (* RS_HS = "m_axi_in_15_R.valid" *)input m_axi_in_15_RVALID;
  (* RS_HS = "m_axi_in_15_W.data" *)output [255:0] m_axi_in_15_WDATA;
  (* RS_HS = "m_axi_in_15_W.data" *)output m_axi_in_15_WLAST;
  (* RS_HS = "m_axi_in_15_W.ready" *)input m_axi_in_15_WREADY;
  (* RS_HS = "m_axi_in_15_W.data" *)output [31:0] m_axi_in_15_WSTRB;
  (* RS_HS = "m_axi_in_15_W.valid" *)output m_axi_in_15_WVALID;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [63:0] m_axi_in_16_ARADDR;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [1:0] m_axi_in_16_ARBURST;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [3:0] m_axi_in_16_ARCACHE;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [0:0] m_axi_in_16_ARID;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [7:0] m_axi_in_16_ARLEN;
  (* RS_HS = "m_axi_in_16_AR.data" *)output m_axi_in_16_ARLOCK;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [2:0] m_axi_in_16_ARPROT;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [3:0] m_axi_in_16_ARQOS;
  (* RS_HS = "m_axi_in_16_AR.ready" *)input m_axi_in_16_ARREADY;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [2:0] m_axi_in_16_ARSIZE;
  (* RS_HS = "m_axi_in_16_AR.valid" *)output m_axi_in_16_ARVALID;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [63:0] m_axi_in_16_AWADDR;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [1:0] m_axi_in_16_AWBURST;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [3:0] m_axi_in_16_AWCACHE;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [0:0] m_axi_in_16_AWID;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [7:0] m_axi_in_16_AWLEN;
  (* RS_HS = "m_axi_in_16_AW.data" *)output m_axi_in_16_AWLOCK;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [2:0] m_axi_in_16_AWPROT;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [3:0] m_axi_in_16_AWQOS;
  (* RS_HS = "m_axi_in_16_AW.ready" *)input m_axi_in_16_AWREADY;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [2:0] m_axi_in_16_AWSIZE;
  (* RS_HS = "m_axi_in_16_AW.valid" *)output m_axi_in_16_AWVALID;
  (* RS_HS = "m_axi_in_16_B.data" *)input [0:0] m_axi_in_16_BID;
  (* RS_HS = "m_axi_in_16_B.ready" *)output m_axi_in_16_BREADY;
  (* RS_HS = "m_axi_in_16_B.data" *)input [1:0] m_axi_in_16_BRESP;
  (* RS_HS = "m_axi_in_16_B.valid" *)input m_axi_in_16_BVALID;
  (* RS_HS = "m_axi_in_16_R.data" *)input [255:0] m_axi_in_16_RDATA;
  (* RS_HS = "m_axi_in_16_R.data" *)input [0:0] m_axi_in_16_RID;
  (* RS_HS = "m_axi_in_16_R.data" *)input m_axi_in_16_RLAST;
  (* RS_HS = "m_axi_in_16_R.ready" *)output m_axi_in_16_RREADY;
  (* RS_HS = "m_axi_in_16_R.data" *)input [1:0] m_axi_in_16_RRESP;
  (* RS_HS = "m_axi_in_16_R.valid" *)input m_axi_in_16_RVALID;
  (* RS_HS = "m_axi_in_16_W.data" *)output [255:0] m_axi_in_16_WDATA;
  (* RS_HS = "m_axi_in_16_W.data" *)output m_axi_in_16_WLAST;
  (* RS_HS = "m_axi_in_16_W.ready" *)input m_axi_in_16_WREADY;
  (* RS_HS = "m_axi_in_16_W.data" *)output [31:0] m_axi_in_16_WSTRB;
  (* RS_HS = "m_axi_in_16_W.valid" *)output m_axi_in_16_WVALID;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [63:0] m_axi_in_17_ARADDR;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [1:0] m_axi_in_17_ARBURST;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [3:0] m_axi_in_17_ARCACHE;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [0:0] m_axi_in_17_ARID;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [7:0] m_axi_in_17_ARLEN;
  (* RS_HS = "m_axi_in_17_AR.data" *)output m_axi_in_17_ARLOCK;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [2:0] m_axi_in_17_ARPROT;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [3:0] m_axi_in_17_ARQOS;
  (* RS_HS = "m_axi_in_17_AR.ready" *)input m_axi_in_17_ARREADY;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [2:0] m_axi_in_17_ARSIZE;
  (* RS_HS = "m_axi_in_17_AR.valid" *)output m_axi_in_17_ARVALID;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [63:0] m_axi_in_17_AWADDR;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [1:0] m_axi_in_17_AWBURST;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [3:0] m_axi_in_17_AWCACHE;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [0:0] m_axi_in_17_AWID;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [7:0] m_axi_in_17_AWLEN;
  (* RS_HS = "m_axi_in_17_AW.data" *)output m_axi_in_17_AWLOCK;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [2:0] m_axi_in_17_AWPROT;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [3:0] m_axi_in_17_AWQOS;
  (* RS_HS = "m_axi_in_17_AW.ready" *)input m_axi_in_17_AWREADY;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [2:0] m_axi_in_17_AWSIZE;
  (* RS_HS = "m_axi_in_17_AW.valid" *)output m_axi_in_17_AWVALID;
  (* RS_HS = "m_axi_in_17_B.data" *)input [0:0] m_axi_in_17_BID;
  (* RS_HS = "m_axi_in_17_B.ready" *)output m_axi_in_17_BREADY;
  (* RS_HS = "m_axi_in_17_B.data" *)input [1:0] m_axi_in_17_BRESP;
  (* RS_HS = "m_axi_in_17_B.valid" *)input m_axi_in_17_BVALID;
  (* RS_HS = "m_axi_in_17_R.data" *)input [255:0] m_axi_in_17_RDATA;
  (* RS_HS = "m_axi_in_17_R.data" *)input [0:0] m_axi_in_17_RID;
  (* RS_HS = "m_axi_in_17_R.data" *)input m_axi_in_17_RLAST;
  (* RS_HS = "m_axi_in_17_R.ready" *)output m_axi_in_17_RREADY;
  (* RS_HS = "m_axi_in_17_R.data" *)input [1:0] m_axi_in_17_RRESP;
  (* RS_HS = "m_axi_in_17_R.valid" *)input m_axi_in_17_RVALID;
  (* RS_HS = "m_axi_in_17_W.data" *)output [255:0] m_axi_in_17_WDATA;
  (* RS_HS = "m_axi_in_17_W.data" *)output m_axi_in_17_WLAST;
  (* RS_HS = "m_axi_in_17_W.ready" *)input m_axi_in_17_WREADY;
  (* RS_HS = "m_axi_in_17_W.data" *)output [31:0] m_axi_in_17_WSTRB;
  (* RS_HS = "m_axi_in_17_W.valid" *)output m_axi_in_17_WVALID;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [63:0] m_axi_in_18_ARADDR;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [1:0] m_axi_in_18_ARBURST;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [3:0] m_axi_in_18_ARCACHE;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [0:0] m_axi_in_18_ARID;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [7:0] m_axi_in_18_ARLEN;
  (* RS_HS = "m_axi_in_18_AR.data" *)output m_axi_in_18_ARLOCK;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [2:0] m_axi_in_18_ARPROT;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [3:0] m_axi_in_18_ARQOS;
  (* RS_HS = "m_axi_in_18_AR.ready" *)input m_axi_in_18_ARREADY;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [2:0] m_axi_in_18_ARSIZE;
  (* RS_HS = "m_axi_in_18_AR.valid" *)output m_axi_in_18_ARVALID;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [63:0] m_axi_in_18_AWADDR;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [1:0] m_axi_in_18_AWBURST;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [3:0] m_axi_in_18_AWCACHE;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [0:0] m_axi_in_18_AWID;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [7:0] m_axi_in_18_AWLEN;
  (* RS_HS = "m_axi_in_18_AW.data" *)output m_axi_in_18_AWLOCK;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [2:0] m_axi_in_18_AWPROT;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [3:0] m_axi_in_18_AWQOS;
  (* RS_HS = "m_axi_in_18_AW.ready" *)input m_axi_in_18_AWREADY;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [2:0] m_axi_in_18_AWSIZE;
  (* RS_HS = "m_axi_in_18_AW.valid" *)output m_axi_in_18_AWVALID;
  (* RS_HS = "m_axi_in_18_B.data" *)input [0:0] m_axi_in_18_BID;
  (* RS_HS = "m_axi_in_18_B.ready" *)output m_axi_in_18_BREADY;
  (* RS_HS = "m_axi_in_18_B.data" *)input [1:0] m_axi_in_18_BRESP;
  (* RS_HS = "m_axi_in_18_B.valid" *)input m_axi_in_18_BVALID;
  (* RS_HS = "m_axi_in_18_R.data" *)input [255:0] m_axi_in_18_RDATA;
  (* RS_HS = "m_axi_in_18_R.data" *)input [0:0] m_axi_in_18_RID;
  (* RS_HS = "m_axi_in_18_R.data" *)input m_axi_in_18_RLAST;
  (* RS_HS = "m_axi_in_18_R.ready" *)output m_axi_in_18_RREADY;
  (* RS_HS = "m_axi_in_18_R.data" *)input [1:0] m_axi_in_18_RRESP;
  (* RS_HS = "m_axi_in_18_R.valid" *)input m_axi_in_18_RVALID;
  (* RS_HS = "m_axi_in_18_W.data" *)output [255:0] m_axi_in_18_WDATA;
  (* RS_HS = "m_axi_in_18_W.data" *)output m_axi_in_18_WLAST;
  (* RS_HS = "m_axi_in_18_W.ready" *)input m_axi_in_18_WREADY;
  (* RS_HS = "m_axi_in_18_W.data" *)output [31:0] m_axi_in_18_WSTRB;
  (* RS_HS = "m_axi_in_18_W.valid" *)output m_axi_in_18_WVALID;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [63:0] m_axi_in_19_ARADDR;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [1:0] m_axi_in_19_ARBURST;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [3:0] m_axi_in_19_ARCACHE;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [0:0] m_axi_in_19_ARID;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [7:0] m_axi_in_19_ARLEN;
  (* RS_HS = "m_axi_in_19_AR.data" *)output m_axi_in_19_ARLOCK;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [2:0] m_axi_in_19_ARPROT;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [3:0] m_axi_in_19_ARQOS;
  (* RS_HS = "m_axi_in_19_AR.ready" *)input m_axi_in_19_ARREADY;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [2:0] m_axi_in_19_ARSIZE;
  (* RS_HS = "m_axi_in_19_AR.valid" *)output m_axi_in_19_ARVALID;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [63:0] m_axi_in_19_AWADDR;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [1:0] m_axi_in_19_AWBURST;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [3:0] m_axi_in_19_AWCACHE;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [0:0] m_axi_in_19_AWID;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [7:0] m_axi_in_19_AWLEN;
  (* RS_HS = "m_axi_in_19_AW.data" *)output m_axi_in_19_AWLOCK;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [2:0] m_axi_in_19_AWPROT;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [3:0] m_axi_in_19_AWQOS;
  (* RS_HS = "m_axi_in_19_AW.ready" *)input m_axi_in_19_AWREADY;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [2:0] m_axi_in_19_AWSIZE;
  (* RS_HS = "m_axi_in_19_AW.valid" *)output m_axi_in_19_AWVALID;
  (* RS_HS = "m_axi_in_19_B.data" *)input [0:0] m_axi_in_19_BID;
  (* RS_HS = "m_axi_in_19_B.ready" *)output m_axi_in_19_BREADY;
  (* RS_HS = "m_axi_in_19_B.data" *)input [1:0] m_axi_in_19_BRESP;
  (* RS_HS = "m_axi_in_19_B.valid" *)input m_axi_in_19_BVALID;
  (* RS_HS = "m_axi_in_19_R.data" *)input [255:0] m_axi_in_19_RDATA;
  (* RS_HS = "m_axi_in_19_R.data" *)input [0:0] m_axi_in_19_RID;
  (* RS_HS = "m_axi_in_19_R.data" *)input m_axi_in_19_RLAST;
  (* RS_HS = "m_axi_in_19_R.ready" *)output m_axi_in_19_RREADY;
  (* RS_HS = "m_axi_in_19_R.data" *)input [1:0] m_axi_in_19_RRESP;
  (* RS_HS = "m_axi_in_19_R.valid" *)input m_axi_in_19_RVALID;
  (* RS_HS = "m_axi_in_19_W.data" *)output [255:0] m_axi_in_19_WDATA;
  (* RS_HS = "m_axi_in_19_W.data" *)output m_axi_in_19_WLAST;
  (* RS_HS = "m_axi_in_19_W.ready" *)input m_axi_in_19_WREADY;
  (* RS_HS = "m_axi_in_19_W.data" *)output [31:0] m_axi_in_19_WSTRB;
  (* RS_HS = "m_axi_in_19_W.valid" *)output m_axi_in_19_WVALID;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [63:0] m_axi_in_2_ARADDR;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [1:0] m_axi_in_2_ARBURST;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [3:0] m_axi_in_2_ARCACHE;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [0:0] m_axi_in_2_ARID;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [7:0] m_axi_in_2_ARLEN;
  (* RS_HS = "m_axi_in_2_AR.data" *)output m_axi_in_2_ARLOCK;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [2:0] m_axi_in_2_ARPROT;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [3:0] m_axi_in_2_ARQOS;
  (* RS_HS = "m_axi_in_2_AR.ready" *)input m_axi_in_2_ARREADY;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [2:0] m_axi_in_2_ARSIZE;
  (* RS_HS = "m_axi_in_2_AR.valid" *)output m_axi_in_2_ARVALID;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [63:0] m_axi_in_2_AWADDR;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [1:0] m_axi_in_2_AWBURST;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [3:0] m_axi_in_2_AWCACHE;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [0:0] m_axi_in_2_AWID;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [7:0] m_axi_in_2_AWLEN;
  (* RS_HS = "m_axi_in_2_AW.data" *)output m_axi_in_2_AWLOCK;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [2:0] m_axi_in_2_AWPROT;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [3:0] m_axi_in_2_AWQOS;
  (* RS_HS = "m_axi_in_2_AW.ready" *)input m_axi_in_2_AWREADY;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [2:0] m_axi_in_2_AWSIZE;
  (* RS_HS = "m_axi_in_2_AW.valid" *)output m_axi_in_2_AWVALID;
  (* RS_HS = "m_axi_in_2_B.data" *)input [0:0] m_axi_in_2_BID;
  (* RS_HS = "m_axi_in_2_B.ready" *)output m_axi_in_2_BREADY;
  (* RS_HS = "m_axi_in_2_B.data" *)input [1:0] m_axi_in_2_BRESP;
  (* RS_HS = "m_axi_in_2_B.valid" *)input m_axi_in_2_BVALID;
  (* RS_HS = "m_axi_in_2_R.data" *)input [255:0] m_axi_in_2_RDATA;
  (* RS_HS = "m_axi_in_2_R.data" *)input [0:0] m_axi_in_2_RID;
  (* RS_HS = "m_axi_in_2_R.data" *)input m_axi_in_2_RLAST;
  (* RS_HS = "m_axi_in_2_R.ready" *)output m_axi_in_2_RREADY;
  (* RS_HS = "m_axi_in_2_R.data" *)input [1:0] m_axi_in_2_RRESP;
  (* RS_HS = "m_axi_in_2_R.valid" *)input m_axi_in_2_RVALID;
  (* RS_HS = "m_axi_in_2_W.data" *)output [255:0] m_axi_in_2_WDATA;
  (* RS_HS = "m_axi_in_2_W.data" *)output m_axi_in_2_WLAST;
  (* RS_HS = "m_axi_in_2_W.ready" *)input m_axi_in_2_WREADY;
  (* RS_HS = "m_axi_in_2_W.data" *)output [31:0] m_axi_in_2_WSTRB;
  (* RS_HS = "m_axi_in_2_W.valid" *)output m_axi_in_2_WVALID;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [63:0] m_axi_in_20_ARADDR;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [1:0] m_axi_in_20_ARBURST;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [3:0] m_axi_in_20_ARCACHE;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [0:0] m_axi_in_20_ARID;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [7:0] m_axi_in_20_ARLEN;
  (* RS_HS = "m_axi_in_20_AR.data" *)output m_axi_in_20_ARLOCK;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [2:0] m_axi_in_20_ARPROT;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [3:0] m_axi_in_20_ARQOS;
  (* RS_HS = "m_axi_in_20_AR.ready" *)input m_axi_in_20_ARREADY;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [2:0] m_axi_in_20_ARSIZE;
  (* RS_HS = "m_axi_in_20_AR.valid" *)output m_axi_in_20_ARVALID;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [63:0] m_axi_in_20_AWADDR;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [1:0] m_axi_in_20_AWBURST;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [3:0] m_axi_in_20_AWCACHE;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [0:0] m_axi_in_20_AWID;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [7:0] m_axi_in_20_AWLEN;
  (* RS_HS = "m_axi_in_20_AW.data" *)output m_axi_in_20_AWLOCK;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [2:0] m_axi_in_20_AWPROT;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [3:0] m_axi_in_20_AWQOS;
  (* RS_HS = "m_axi_in_20_AW.ready" *)input m_axi_in_20_AWREADY;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [2:0] m_axi_in_20_AWSIZE;
  (* RS_HS = "m_axi_in_20_AW.valid" *)output m_axi_in_20_AWVALID;
  (* RS_HS = "m_axi_in_20_B.data" *)input [0:0] m_axi_in_20_BID;
  (* RS_HS = "m_axi_in_20_B.ready" *)output m_axi_in_20_BREADY;
  (* RS_HS = "m_axi_in_20_B.data" *)input [1:0] m_axi_in_20_BRESP;
  (* RS_HS = "m_axi_in_20_B.valid" *)input m_axi_in_20_BVALID;
  (* RS_HS = "m_axi_in_20_R.data" *)input [255:0] m_axi_in_20_RDATA;
  (* RS_HS = "m_axi_in_20_R.data" *)input [0:0] m_axi_in_20_RID;
  (* RS_HS = "m_axi_in_20_R.data" *)input m_axi_in_20_RLAST;
  (* RS_HS = "m_axi_in_20_R.ready" *)output m_axi_in_20_RREADY;
  (* RS_HS = "m_axi_in_20_R.data" *)input [1:0] m_axi_in_20_RRESP;
  (* RS_HS = "m_axi_in_20_R.valid" *)input m_axi_in_20_RVALID;
  (* RS_HS = "m_axi_in_20_W.data" *)output [255:0] m_axi_in_20_WDATA;
  (* RS_HS = "m_axi_in_20_W.data" *)output m_axi_in_20_WLAST;
  (* RS_HS = "m_axi_in_20_W.ready" *)input m_axi_in_20_WREADY;
  (* RS_HS = "m_axi_in_20_W.data" *)output [31:0] m_axi_in_20_WSTRB;
  (* RS_HS = "m_axi_in_20_W.valid" *)output m_axi_in_20_WVALID;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [63:0] m_axi_in_21_ARADDR;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [1:0] m_axi_in_21_ARBURST;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [3:0] m_axi_in_21_ARCACHE;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [0:0] m_axi_in_21_ARID;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [7:0] m_axi_in_21_ARLEN;
  (* RS_HS = "m_axi_in_21_AR.data" *)output m_axi_in_21_ARLOCK;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [2:0] m_axi_in_21_ARPROT;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [3:0] m_axi_in_21_ARQOS;
  (* RS_HS = "m_axi_in_21_AR.ready" *)input m_axi_in_21_ARREADY;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [2:0] m_axi_in_21_ARSIZE;
  (* RS_HS = "m_axi_in_21_AR.valid" *)output m_axi_in_21_ARVALID;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [63:0] m_axi_in_21_AWADDR;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [1:0] m_axi_in_21_AWBURST;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [3:0] m_axi_in_21_AWCACHE;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [0:0] m_axi_in_21_AWID;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [7:0] m_axi_in_21_AWLEN;
  (* RS_HS = "m_axi_in_21_AW.data" *)output m_axi_in_21_AWLOCK;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [2:0] m_axi_in_21_AWPROT;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [3:0] m_axi_in_21_AWQOS;
  (* RS_HS = "m_axi_in_21_AW.ready" *)input m_axi_in_21_AWREADY;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [2:0] m_axi_in_21_AWSIZE;
  (* RS_HS = "m_axi_in_21_AW.valid" *)output m_axi_in_21_AWVALID;
  (* RS_HS = "m_axi_in_21_B.data" *)input [0:0] m_axi_in_21_BID;
  (* RS_HS = "m_axi_in_21_B.ready" *)output m_axi_in_21_BREADY;
  (* RS_HS = "m_axi_in_21_B.data" *)input [1:0] m_axi_in_21_BRESP;
  (* RS_HS = "m_axi_in_21_B.valid" *)input m_axi_in_21_BVALID;
  (* RS_HS = "m_axi_in_21_R.data" *)input [255:0] m_axi_in_21_RDATA;
  (* RS_HS = "m_axi_in_21_R.data" *)input [0:0] m_axi_in_21_RID;
  (* RS_HS = "m_axi_in_21_R.data" *)input m_axi_in_21_RLAST;
  (* RS_HS = "m_axi_in_21_R.ready" *)output m_axi_in_21_RREADY;
  (* RS_HS = "m_axi_in_21_R.data" *)input [1:0] m_axi_in_21_RRESP;
  (* RS_HS = "m_axi_in_21_R.valid" *)input m_axi_in_21_RVALID;
  (* RS_HS = "m_axi_in_21_W.data" *)output [255:0] m_axi_in_21_WDATA;
  (* RS_HS = "m_axi_in_21_W.data" *)output m_axi_in_21_WLAST;
  (* RS_HS = "m_axi_in_21_W.ready" *)input m_axi_in_21_WREADY;
  (* RS_HS = "m_axi_in_21_W.data" *)output [31:0] m_axi_in_21_WSTRB;
  (* RS_HS = "m_axi_in_21_W.valid" *)output m_axi_in_21_WVALID;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [63:0] m_axi_in_22_ARADDR;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [1:0] m_axi_in_22_ARBURST;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [3:0] m_axi_in_22_ARCACHE;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [0:0] m_axi_in_22_ARID;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [7:0] m_axi_in_22_ARLEN;
  (* RS_HS = "m_axi_in_22_AR.data" *)output m_axi_in_22_ARLOCK;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [2:0] m_axi_in_22_ARPROT;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [3:0] m_axi_in_22_ARQOS;
  (* RS_HS = "m_axi_in_22_AR.ready" *)input m_axi_in_22_ARREADY;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [2:0] m_axi_in_22_ARSIZE;
  (* RS_HS = "m_axi_in_22_AR.valid" *)output m_axi_in_22_ARVALID;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [63:0] m_axi_in_22_AWADDR;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [1:0] m_axi_in_22_AWBURST;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [3:0] m_axi_in_22_AWCACHE;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [0:0] m_axi_in_22_AWID;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [7:0] m_axi_in_22_AWLEN;
  (* RS_HS = "m_axi_in_22_AW.data" *)output m_axi_in_22_AWLOCK;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [2:0] m_axi_in_22_AWPROT;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [3:0] m_axi_in_22_AWQOS;
  (* RS_HS = "m_axi_in_22_AW.ready" *)input m_axi_in_22_AWREADY;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [2:0] m_axi_in_22_AWSIZE;
  (* RS_HS = "m_axi_in_22_AW.valid" *)output m_axi_in_22_AWVALID;
  (* RS_HS = "m_axi_in_22_B.data" *)input [0:0] m_axi_in_22_BID;
  (* RS_HS = "m_axi_in_22_B.ready" *)output m_axi_in_22_BREADY;
  (* RS_HS = "m_axi_in_22_B.data" *)input [1:0] m_axi_in_22_BRESP;
  (* RS_HS = "m_axi_in_22_B.valid" *)input m_axi_in_22_BVALID;
  (* RS_HS = "m_axi_in_22_R.data" *)input [255:0] m_axi_in_22_RDATA;
  (* RS_HS = "m_axi_in_22_R.data" *)input [0:0] m_axi_in_22_RID;
  (* RS_HS = "m_axi_in_22_R.data" *)input m_axi_in_22_RLAST;
  (* RS_HS = "m_axi_in_22_R.ready" *)output m_axi_in_22_RREADY;
  (* RS_HS = "m_axi_in_22_R.data" *)input [1:0] m_axi_in_22_RRESP;
  (* RS_HS = "m_axi_in_22_R.valid" *)input m_axi_in_22_RVALID;
  (* RS_HS = "m_axi_in_22_W.data" *)output [255:0] m_axi_in_22_WDATA;
  (* RS_HS = "m_axi_in_22_W.data" *)output m_axi_in_22_WLAST;
  (* RS_HS = "m_axi_in_22_W.ready" *)input m_axi_in_22_WREADY;
  (* RS_HS = "m_axi_in_22_W.data" *)output [31:0] m_axi_in_22_WSTRB;
  (* RS_HS = "m_axi_in_22_W.valid" *)output m_axi_in_22_WVALID;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [63:0] m_axi_in_23_ARADDR;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [1:0] m_axi_in_23_ARBURST;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [3:0] m_axi_in_23_ARCACHE;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [0:0] m_axi_in_23_ARID;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [7:0] m_axi_in_23_ARLEN;
  (* RS_HS = "m_axi_in_23_AR.data" *)output m_axi_in_23_ARLOCK;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [2:0] m_axi_in_23_ARPROT;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [3:0] m_axi_in_23_ARQOS;
  (* RS_HS = "m_axi_in_23_AR.ready" *)input m_axi_in_23_ARREADY;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [2:0] m_axi_in_23_ARSIZE;
  (* RS_HS = "m_axi_in_23_AR.valid" *)output m_axi_in_23_ARVALID;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [63:0] m_axi_in_23_AWADDR;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [1:0] m_axi_in_23_AWBURST;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [3:0] m_axi_in_23_AWCACHE;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [0:0] m_axi_in_23_AWID;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [7:0] m_axi_in_23_AWLEN;
  (* RS_HS = "m_axi_in_23_AW.data" *)output m_axi_in_23_AWLOCK;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [2:0] m_axi_in_23_AWPROT;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [3:0] m_axi_in_23_AWQOS;
  (* RS_HS = "m_axi_in_23_AW.ready" *)input m_axi_in_23_AWREADY;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [2:0] m_axi_in_23_AWSIZE;
  (* RS_HS = "m_axi_in_23_AW.valid" *)output m_axi_in_23_AWVALID;
  (* RS_HS = "m_axi_in_23_B.data" *)input [0:0] m_axi_in_23_BID;
  (* RS_HS = "m_axi_in_23_B.ready" *)output m_axi_in_23_BREADY;
  (* RS_HS = "m_axi_in_23_B.data" *)input [1:0] m_axi_in_23_BRESP;
  (* RS_HS = "m_axi_in_23_B.valid" *)input m_axi_in_23_BVALID;
  (* RS_HS = "m_axi_in_23_R.data" *)input [255:0] m_axi_in_23_RDATA;
  (* RS_HS = "m_axi_in_23_R.data" *)input [0:0] m_axi_in_23_RID;
  (* RS_HS = "m_axi_in_23_R.data" *)input m_axi_in_23_RLAST;
  (* RS_HS = "m_axi_in_23_R.ready" *)output m_axi_in_23_RREADY;
  (* RS_HS = "m_axi_in_23_R.data" *)input [1:0] m_axi_in_23_RRESP;
  (* RS_HS = "m_axi_in_23_R.valid" *)input m_axi_in_23_RVALID;
  (* RS_HS = "m_axi_in_23_W.data" *)output [255:0] m_axi_in_23_WDATA;
  (* RS_HS = "m_axi_in_23_W.data" *)output m_axi_in_23_WLAST;
  (* RS_HS = "m_axi_in_23_W.ready" *)input m_axi_in_23_WREADY;
  (* RS_HS = "m_axi_in_23_W.data" *)output [31:0] m_axi_in_23_WSTRB;
  (* RS_HS = "m_axi_in_23_W.valid" *)output m_axi_in_23_WVALID;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [63:0] m_axi_in_24_ARADDR;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [1:0] m_axi_in_24_ARBURST;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [3:0] m_axi_in_24_ARCACHE;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [0:0] m_axi_in_24_ARID;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [7:0] m_axi_in_24_ARLEN;
  (* RS_HS = "m_axi_in_24_AR.data" *)output m_axi_in_24_ARLOCK;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [2:0] m_axi_in_24_ARPROT;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [3:0] m_axi_in_24_ARQOS;
  (* RS_HS = "m_axi_in_24_AR.ready" *)input m_axi_in_24_ARREADY;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [2:0] m_axi_in_24_ARSIZE;
  (* RS_HS = "m_axi_in_24_AR.valid" *)output m_axi_in_24_ARVALID;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [63:0] m_axi_in_24_AWADDR;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [1:0] m_axi_in_24_AWBURST;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [3:0] m_axi_in_24_AWCACHE;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [0:0] m_axi_in_24_AWID;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [7:0] m_axi_in_24_AWLEN;
  (* RS_HS = "m_axi_in_24_AW.data" *)output m_axi_in_24_AWLOCK;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [2:0] m_axi_in_24_AWPROT;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [3:0] m_axi_in_24_AWQOS;
  (* RS_HS = "m_axi_in_24_AW.ready" *)input m_axi_in_24_AWREADY;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [2:0] m_axi_in_24_AWSIZE;
  (* RS_HS = "m_axi_in_24_AW.valid" *)output m_axi_in_24_AWVALID;
  (* RS_HS = "m_axi_in_24_B.data" *)input [0:0] m_axi_in_24_BID;
  (* RS_HS = "m_axi_in_24_B.ready" *)output m_axi_in_24_BREADY;
  (* RS_HS = "m_axi_in_24_B.data" *)input [1:0] m_axi_in_24_BRESP;
  (* RS_HS = "m_axi_in_24_B.valid" *)input m_axi_in_24_BVALID;
  (* RS_HS = "m_axi_in_24_R.data" *)input [255:0] m_axi_in_24_RDATA;
  (* RS_HS = "m_axi_in_24_R.data" *)input [0:0] m_axi_in_24_RID;
  (* RS_HS = "m_axi_in_24_R.data" *)input m_axi_in_24_RLAST;
  (* RS_HS = "m_axi_in_24_R.ready" *)output m_axi_in_24_RREADY;
  (* RS_HS = "m_axi_in_24_R.data" *)input [1:0] m_axi_in_24_RRESP;
  (* RS_HS = "m_axi_in_24_R.valid" *)input m_axi_in_24_RVALID;
  (* RS_HS = "m_axi_in_24_W.data" *)output [255:0] m_axi_in_24_WDATA;
  (* RS_HS = "m_axi_in_24_W.data" *)output m_axi_in_24_WLAST;
  (* RS_HS = "m_axi_in_24_W.ready" *)input m_axi_in_24_WREADY;
  (* RS_HS = "m_axi_in_24_W.data" *)output [31:0] m_axi_in_24_WSTRB;
  (* RS_HS = "m_axi_in_24_W.valid" *)output m_axi_in_24_WVALID;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [63:0] m_axi_in_25_ARADDR;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [1:0] m_axi_in_25_ARBURST;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [3:0] m_axi_in_25_ARCACHE;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [0:0] m_axi_in_25_ARID;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [7:0] m_axi_in_25_ARLEN;
  (* RS_HS = "m_axi_in_25_AR.data" *)output m_axi_in_25_ARLOCK;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [2:0] m_axi_in_25_ARPROT;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [3:0] m_axi_in_25_ARQOS;
  (* RS_HS = "m_axi_in_25_AR.ready" *)input m_axi_in_25_ARREADY;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [2:0] m_axi_in_25_ARSIZE;
  (* RS_HS = "m_axi_in_25_AR.valid" *)output m_axi_in_25_ARVALID;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [63:0] m_axi_in_25_AWADDR;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [1:0] m_axi_in_25_AWBURST;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [3:0] m_axi_in_25_AWCACHE;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [0:0] m_axi_in_25_AWID;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [7:0] m_axi_in_25_AWLEN;
  (* RS_HS = "m_axi_in_25_AW.data" *)output m_axi_in_25_AWLOCK;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [2:0] m_axi_in_25_AWPROT;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [3:0] m_axi_in_25_AWQOS;
  (* RS_HS = "m_axi_in_25_AW.ready" *)input m_axi_in_25_AWREADY;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [2:0] m_axi_in_25_AWSIZE;
  (* RS_HS = "m_axi_in_25_AW.valid" *)output m_axi_in_25_AWVALID;
  (* RS_HS = "m_axi_in_25_B.data" *)input [0:0] m_axi_in_25_BID;
  (* RS_HS = "m_axi_in_25_B.ready" *)output m_axi_in_25_BREADY;
  (* RS_HS = "m_axi_in_25_B.data" *)input [1:0] m_axi_in_25_BRESP;
  (* RS_HS = "m_axi_in_25_B.valid" *)input m_axi_in_25_BVALID;
  (* RS_HS = "m_axi_in_25_R.data" *)input [255:0] m_axi_in_25_RDATA;
  (* RS_HS = "m_axi_in_25_R.data" *)input [0:0] m_axi_in_25_RID;
  (* RS_HS = "m_axi_in_25_R.data" *)input m_axi_in_25_RLAST;
  (* RS_HS = "m_axi_in_25_R.ready" *)output m_axi_in_25_RREADY;
  (* RS_HS = "m_axi_in_25_R.data" *)input [1:0] m_axi_in_25_RRESP;
  (* RS_HS = "m_axi_in_25_R.valid" *)input m_axi_in_25_RVALID;
  (* RS_HS = "m_axi_in_25_W.data" *)output [255:0] m_axi_in_25_WDATA;
  (* RS_HS = "m_axi_in_25_W.data" *)output m_axi_in_25_WLAST;
  (* RS_HS = "m_axi_in_25_W.ready" *)input m_axi_in_25_WREADY;
  (* RS_HS = "m_axi_in_25_W.data" *)output [31:0] m_axi_in_25_WSTRB;
  (* RS_HS = "m_axi_in_25_W.valid" *)output m_axi_in_25_WVALID;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [63:0] m_axi_in_26_ARADDR;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [1:0] m_axi_in_26_ARBURST;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [3:0] m_axi_in_26_ARCACHE;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [0:0] m_axi_in_26_ARID;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [7:0] m_axi_in_26_ARLEN;
  (* RS_HS = "m_axi_in_26_AR.data" *)output m_axi_in_26_ARLOCK;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [2:0] m_axi_in_26_ARPROT;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [3:0] m_axi_in_26_ARQOS;
  (* RS_HS = "m_axi_in_26_AR.ready" *)input m_axi_in_26_ARREADY;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [2:0] m_axi_in_26_ARSIZE;
  (* RS_HS = "m_axi_in_26_AR.valid" *)output m_axi_in_26_ARVALID;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [63:0] m_axi_in_26_AWADDR;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [1:0] m_axi_in_26_AWBURST;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [3:0] m_axi_in_26_AWCACHE;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [0:0] m_axi_in_26_AWID;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [7:0] m_axi_in_26_AWLEN;
  (* RS_HS = "m_axi_in_26_AW.data" *)output m_axi_in_26_AWLOCK;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [2:0] m_axi_in_26_AWPROT;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [3:0] m_axi_in_26_AWQOS;
  (* RS_HS = "m_axi_in_26_AW.ready" *)input m_axi_in_26_AWREADY;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [2:0] m_axi_in_26_AWSIZE;
  (* RS_HS = "m_axi_in_26_AW.valid" *)output m_axi_in_26_AWVALID;
  (* RS_HS = "m_axi_in_26_B.data" *)input [0:0] m_axi_in_26_BID;
  (* RS_HS = "m_axi_in_26_B.ready" *)output m_axi_in_26_BREADY;
  (* RS_HS = "m_axi_in_26_B.data" *)input [1:0] m_axi_in_26_BRESP;
  (* RS_HS = "m_axi_in_26_B.valid" *)input m_axi_in_26_BVALID;
  (* RS_HS = "m_axi_in_26_R.data" *)input [255:0] m_axi_in_26_RDATA;
  (* RS_HS = "m_axi_in_26_R.data" *)input [0:0] m_axi_in_26_RID;
  (* RS_HS = "m_axi_in_26_R.data" *)input m_axi_in_26_RLAST;
  (* RS_HS = "m_axi_in_26_R.ready" *)output m_axi_in_26_RREADY;
  (* RS_HS = "m_axi_in_26_R.data" *)input [1:0] m_axi_in_26_RRESP;
  (* RS_HS = "m_axi_in_26_R.valid" *)input m_axi_in_26_RVALID;
  (* RS_HS = "m_axi_in_26_W.data" *)output [255:0] m_axi_in_26_WDATA;
  (* RS_HS = "m_axi_in_26_W.data" *)output m_axi_in_26_WLAST;
  (* RS_HS = "m_axi_in_26_W.ready" *)input m_axi_in_26_WREADY;
  (* RS_HS = "m_axi_in_26_W.data" *)output [31:0] m_axi_in_26_WSTRB;
  (* RS_HS = "m_axi_in_26_W.valid" *)output m_axi_in_26_WVALID;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [63:0] m_axi_in_27_ARADDR;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [1:0] m_axi_in_27_ARBURST;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [3:0] m_axi_in_27_ARCACHE;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [0:0] m_axi_in_27_ARID;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [7:0] m_axi_in_27_ARLEN;
  (* RS_HS = "m_axi_in_27_AR.data" *)output m_axi_in_27_ARLOCK;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [2:0] m_axi_in_27_ARPROT;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [3:0] m_axi_in_27_ARQOS;
  (* RS_HS = "m_axi_in_27_AR.ready" *)input m_axi_in_27_ARREADY;
  (* RS_HS = "m_axi_in_27_AR.data" *)output [2:0] m_axi_in_27_ARSIZE;
  (* RS_HS = "m_axi_in_27_AR.valid" *)output m_axi_in_27_ARVALID;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [63:0] m_axi_in_27_AWADDR;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [1:0] m_axi_in_27_AWBURST;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [3:0] m_axi_in_27_AWCACHE;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [0:0] m_axi_in_27_AWID;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [7:0] m_axi_in_27_AWLEN;
  (* RS_HS = "m_axi_in_27_AW.data" *)output m_axi_in_27_AWLOCK;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [2:0] m_axi_in_27_AWPROT;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [3:0] m_axi_in_27_AWQOS;
  (* RS_HS = "m_axi_in_27_AW.ready" *)input m_axi_in_27_AWREADY;
  (* RS_HS = "m_axi_in_27_AW.data" *)output [2:0] m_axi_in_27_AWSIZE;
  (* RS_HS = "m_axi_in_27_AW.valid" *)output m_axi_in_27_AWVALID;
  (* RS_HS = "m_axi_in_27_B.data" *)input [0:0] m_axi_in_27_BID;
  (* RS_HS = "m_axi_in_27_B.ready" *)output m_axi_in_27_BREADY;
  (* RS_HS = "m_axi_in_27_B.data" *)input [1:0] m_axi_in_27_BRESP;
  (* RS_HS = "m_axi_in_27_B.valid" *)input m_axi_in_27_BVALID;
  (* RS_HS = "m_axi_in_27_R.data" *)input [255:0] m_axi_in_27_RDATA;
  (* RS_HS = "m_axi_in_27_R.data" *)input [0:0] m_axi_in_27_RID;
  (* RS_HS = "m_axi_in_27_R.data" *)input m_axi_in_27_RLAST;
  (* RS_HS = "m_axi_in_27_R.ready" *)output m_axi_in_27_RREADY;
  (* RS_HS = "m_axi_in_27_R.data" *)input [1:0] m_axi_in_27_RRESP;
  (* RS_HS = "m_axi_in_27_R.valid" *)input m_axi_in_27_RVALID;
  (* RS_HS = "m_axi_in_27_W.data" *)output [255:0] m_axi_in_27_WDATA;
  (* RS_HS = "m_axi_in_27_W.data" *)output m_axi_in_27_WLAST;
  (* RS_HS = "m_axi_in_27_W.ready" *)input m_axi_in_27_WREADY;
  (* RS_HS = "m_axi_in_27_W.data" *)output [31:0] m_axi_in_27_WSTRB;
  (* RS_HS = "m_axi_in_27_W.valid" *)output m_axi_in_27_WVALID;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [63:0] m_axi_in_28_ARADDR;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [1:0] m_axi_in_28_ARBURST;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [3:0] m_axi_in_28_ARCACHE;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [0:0] m_axi_in_28_ARID;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [7:0] m_axi_in_28_ARLEN;
  (* RS_HS = "m_axi_in_28_AR.data" *)output m_axi_in_28_ARLOCK;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [2:0] m_axi_in_28_ARPROT;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [3:0] m_axi_in_28_ARQOS;
  (* RS_HS = "m_axi_in_28_AR.ready" *)input m_axi_in_28_ARREADY;
  (* RS_HS = "m_axi_in_28_AR.data" *)output [2:0] m_axi_in_28_ARSIZE;
  (* RS_HS = "m_axi_in_28_AR.valid" *)output m_axi_in_28_ARVALID;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [63:0] m_axi_in_28_AWADDR;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [1:0] m_axi_in_28_AWBURST;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [3:0] m_axi_in_28_AWCACHE;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [0:0] m_axi_in_28_AWID;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [7:0] m_axi_in_28_AWLEN;
  (* RS_HS = "m_axi_in_28_AW.data" *)output m_axi_in_28_AWLOCK;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [2:0] m_axi_in_28_AWPROT;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [3:0] m_axi_in_28_AWQOS;
  (* RS_HS = "m_axi_in_28_AW.ready" *)input m_axi_in_28_AWREADY;
  (* RS_HS = "m_axi_in_28_AW.data" *)output [2:0] m_axi_in_28_AWSIZE;
  (* RS_HS = "m_axi_in_28_AW.valid" *)output m_axi_in_28_AWVALID;
  (* RS_HS = "m_axi_in_28_B.data" *)input [0:0] m_axi_in_28_BID;
  (* RS_HS = "m_axi_in_28_B.ready" *)output m_axi_in_28_BREADY;
  (* RS_HS = "m_axi_in_28_B.data" *)input [1:0] m_axi_in_28_BRESP;
  (* RS_HS = "m_axi_in_28_B.valid" *)input m_axi_in_28_BVALID;
  (* RS_HS = "m_axi_in_28_R.data" *)input [255:0] m_axi_in_28_RDATA;
  (* RS_HS = "m_axi_in_28_R.data" *)input [0:0] m_axi_in_28_RID;
  (* RS_HS = "m_axi_in_28_R.data" *)input m_axi_in_28_RLAST;
  (* RS_HS = "m_axi_in_28_R.ready" *)output m_axi_in_28_RREADY;
  (* RS_HS = "m_axi_in_28_R.data" *)input [1:0] m_axi_in_28_RRESP;
  (* RS_HS = "m_axi_in_28_R.valid" *)input m_axi_in_28_RVALID;
  (* RS_HS = "m_axi_in_28_W.data" *)output [255:0] m_axi_in_28_WDATA;
  (* RS_HS = "m_axi_in_28_W.data" *)output m_axi_in_28_WLAST;
  (* RS_HS = "m_axi_in_28_W.ready" *)input m_axi_in_28_WREADY;
  (* RS_HS = "m_axi_in_28_W.data" *)output [31:0] m_axi_in_28_WSTRB;
  (* RS_HS = "m_axi_in_28_W.valid" *)output m_axi_in_28_WVALID;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [63:0] m_axi_in_29_ARADDR;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [1:0] m_axi_in_29_ARBURST;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [3:0] m_axi_in_29_ARCACHE;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [0:0] m_axi_in_29_ARID;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [7:0] m_axi_in_29_ARLEN;
  (* RS_HS = "m_axi_in_29_AR.data" *)output m_axi_in_29_ARLOCK;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [2:0] m_axi_in_29_ARPROT;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [3:0] m_axi_in_29_ARQOS;
  (* RS_HS = "m_axi_in_29_AR.ready" *)input m_axi_in_29_ARREADY;
  (* RS_HS = "m_axi_in_29_AR.data" *)output [2:0] m_axi_in_29_ARSIZE;
  (* RS_HS = "m_axi_in_29_AR.valid" *)output m_axi_in_29_ARVALID;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [63:0] m_axi_in_29_AWADDR;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [1:0] m_axi_in_29_AWBURST;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [3:0] m_axi_in_29_AWCACHE;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [0:0] m_axi_in_29_AWID;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [7:0] m_axi_in_29_AWLEN;
  (* RS_HS = "m_axi_in_29_AW.data" *)output m_axi_in_29_AWLOCK;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [2:0] m_axi_in_29_AWPROT;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [3:0] m_axi_in_29_AWQOS;
  (* RS_HS = "m_axi_in_29_AW.ready" *)input m_axi_in_29_AWREADY;
  (* RS_HS = "m_axi_in_29_AW.data" *)output [2:0] m_axi_in_29_AWSIZE;
  (* RS_HS = "m_axi_in_29_AW.valid" *)output m_axi_in_29_AWVALID;
  (* RS_HS = "m_axi_in_29_B.data" *)input [0:0] m_axi_in_29_BID;
  (* RS_HS = "m_axi_in_29_B.ready" *)output m_axi_in_29_BREADY;
  (* RS_HS = "m_axi_in_29_B.data" *)input [1:0] m_axi_in_29_BRESP;
  (* RS_HS = "m_axi_in_29_B.valid" *)input m_axi_in_29_BVALID;
  (* RS_HS = "m_axi_in_29_R.data" *)input [255:0] m_axi_in_29_RDATA;
  (* RS_HS = "m_axi_in_29_R.data" *)input [0:0] m_axi_in_29_RID;
  (* RS_HS = "m_axi_in_29_R.data" *)input m_axi_in_29_RLAST;
  (* RS_HS = "m_axi_in_29_R.ready" *)output m_axi_in_29_RREADY;
  (* RS_HS = "m_axi_in_29_R.data" *)input [1:0] m_axi_in_29_RRESP;
  (* RS_HS = "m_axi_in_29_R.valid" *)input m_axi_in_29_RVALID;
  (* RS_HS = "m_axi_in_29_W.data" *)output [255:0] m_axi_in_29_WDATA;
  (* RS_HS = "m_axi_in_29_W.data" *)output m_axi_in_29_WLAST;
  (* RS_HS = "m_axi_in_29_W.ready" *)input m_axi_in_29_WREADY;
  (* RS_HS = "m_axi_in_29_W.data" *)output [31:0] m_axi_in_29_WSTRB;
  (* RS_HS = "m_axi_in_29_W.valid" *)output m_axi_in_29_WVALID;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [63:0] m_axi_in_3_ARADDR;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [1:0] m_axi_in_3_ARBURST;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [3:0] m_axi_in_3_ARCACHE;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [0:0] m_axi_in_3_ARID;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [7:0] m_axi_in_3_ARLEN;
  (* RS_HS = "m_axi_in_3_AR.data" *)output m_axi_in_3_ARLOCK;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [2:0] m_axi_in_3_ARPROT;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [3:0] m_axi_in_3_ARQOS;
  (* RS_HS = "m_axi_in_3_AR.ready" *)input m_axi_in_3_ARREADY;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [2:0] m_axi_in_3_ARSIZE;
  (* RS_HS = "m_axi_in_3_AR.valid" *)output m_axi_in_3_ARVALID;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [63:0] m_axi_in_3_AWADDR;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [1:0] m_axi_in_3_AWBURST;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [3:0] m_axi_in_3_AWCACHE;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [0:0] m_axi_in_3_AWID;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [7:0] m_axi_in_3_AWLEN;
  (* RS_HS = "m_axi_in_3_AW.data" *)output m_axi_in_3_AWLOCK;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [2:0] m_axi_in_3_AWPROT;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [3:0] m_axi_in_3_AWQOS;
  (* RS_HS = "m_axi_in_3_AW.ready" *)input m_axi_in_3_AWREADY;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [2:0] m_axi_in_3_AWSIZE;
  (* RS_HS = "m_axi_in_3_AW.valid" *)output m_axi_in_3_AWVALID;
  (* RS_HS = "m_axi_in_3_B.data" *)input [0:0] m_axi_in_3_BID;
  (* RS_HS = "m_axi_in_3_B.ready" *)output m_axi_in_3_BREADY;
  (* RS_HS = "m_axi_in_3_B.data" *)input [1:0] m_axi_in_3_BRESP;
  (* RS_HS = "m_axi_in_3_B.valid" *)input m_axi_in_3_BVALID;
  (* RS_HS = "m_axi_in_3_R.data" *)input [255:0] m_axi_in_3_RDATA;
  (* RS_HS = "m_axi_in_3_R.data" *)input [0:0] m_axi_in_3_RID;
  (* RS_HS = "m_axi_in_3_R.data" *)input m_axi_in_3_RLAST;
  (* RS_HS = "m_axi_in_3_R.ready" *)output m_axi_in_3_RREADY;
  (* RS_HS = "m_axi_in_3_R.data" *)input [1:0] m_axi_in_3_RRESP;
  (* RS_HS = "m_axi_in_3_R.valid" *)input m_axi_in_3_RVALID;
  (* RS_HS = "m_axi_in_3_W.data" *)output [255:0] m_axi_in_3_WDATA;
  (* RS_HS = "m_axi_in_3_W.data" *)output m_axi_in_3_WLAST;
  (* RS_HS = "m_axi_in_3_W.ready" *)input m_axi_in_3_WREADY;
  (* RS_HS = "m_axi_in_3_W.data" *)output [31:0] m_axi_in_3_WSTRB;
  (* RS_HS = "m_axi_in_3_W.valid" *)output m_axi_in_3_WVALID;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [63:0] m_axi_in_30_ARADDR;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [1:0] m_axi_in_30_ARBURST;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [3:0] m_axi_in_30_ARCACHE;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [0:0] m_axi_in_30_ARID;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [7:0] m_axi_in_30_ARLEN;
  (* RS_HS = "m_axi_in_30_AR.data" *)output m_axi_in_30_ARLOCK;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [2:0] m_axi_in_30_ARPROT;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [3:0] m_axi_in_30_ARQOS;
  (* RS_HS = "m_axi_in_30_AR.ready" *)input m_axi_in_30_ARREADY;
  (* RS_HS = "m_axi_in_30_AR.data" *)output [2:0] m_axi_in_30_ARSIZE;
  (* RS_HS = "m_axi_in_30_AR.valid" *)output m_axi_in_30_ARVALID;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [63:0] m_axi_in_30_AWADDR;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [1:0] m_axi_in_30_AWBURST;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [3:0] m_axi_in_30_AWCACHE;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [0:0] m_axi_in_30_AWID;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [7:0] m_axi_in_30_AWLEN;
  (* RS_HS = "m_axi_in_30_AW.data" *)output m_axi_in_30_AWLOCK;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [2:0] m_axi_in_30_AWPROT;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [3:0] m_axi_in_30_AWQOS;
  (* RS_HS = "m_axi_in_30_AW.ready" *)input m_axi_in_30_AWREADY;
  (* RS_HS = "m_axi_in_30_AW.data" *)output [2:0] m_axi_in_30_AWSIZE;
  (* RS_HS = "m_axi_in_30_AW.valid" *)output m_axi_in_30_AWVALID;
  (* RS_HS = "m_axi_in_30_B.data" *)input [0:0] m_axi_in_30_BID;
  (* RS_HS = "m_axi_in_30_B.ready" *)output m_axi_in_30_BREADY;
  (* RS_HS = "m_axi_in_30_B.data" *)input [1:0] m_axi_in_30_BRESP;
  (* RS_HS = "m_axi_in_30_B.valid" *)input m_axi_in_30_BVALID;
  (* RS_HS = "m_axi_in_30_R.data" *)input [255:0] m_axi_in_30_RDATA;
  (* RS_HS = "m_axi_in_30_R.data" *)input [0:0] m_axi_in_30_RID;
  (* RS_HS = "m_axi_in_30_R.data" *)input m_axi_in_30_RLAST;
  (* RS_HS = "m_axi_in_30_R.ready" *)output m_axi_in_30_RREADY;
  (* RS_HS = "m_axi_in_30_R.data" *)input [1:0] m_axi_in_30_RRESP;
  (* RS_HS = "m_axi_in_30_R.valid" *)input m_axi_in_30_RVALID;
  (* RS_HS = "m_axi_in_30_W.data" *)output [255:0] m_axi_in_30_WDATA;
  (* RS_HS = "m_axi_in_30_W.data" *)output m_axi_in_30_WLAST;
  (* RS_HS = "m_axi_in_30_W.ready" *)input m_axi_in_30_WREADY;
  (* RS_HS = "m_axi_in_30_W.data" *)output [31:0] m_axi_in_30_WSTRB;
  (* RS_HS = "m_axi_in_30_W.valid" *)output m_axi_in_30_WVALID;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [63:0] m_axi_in_31_ARADDR;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [1:0] m_axi_in_31_ARBURST;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [3:0] m_axi_in_31_ARCACHE;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [0:0] m_axi_in_31_ARID;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [7:0] m_axi_in_31_ARLEN;
  (* RS_HS = "m_axi_in_31_AR.data" *)output m_axi_in_31_ARLOCK;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [2:0] m_axi_in_31_ARPROT;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [3:0] m_axi_in_31_ARQOS;
  (* RS_HS = "m_axi_in_31_AR.ready" *)input m_axi_in_31_ARREADY;
  (* RS_HS = "m_axi_in_31_AR.data" *)output [2:0] m_axi_in_31_ARSIZE;
  (* RS_HS = "m_axi_in_31_AR.valid" *)output m_axi_in_31_ARVALID;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [63:0] m_axi_in_31_AWADDR;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [1:0] m_axi_in_31_AWBURST;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [3:0] m_axi_in_31_AWCACHE;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [0:0] m_axi_in_31_AWID;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [7:0] m_axi_in_31_AWLEN;
  (* RS_HS = "m_axi_in_31_AW.data" *)output m_axi_in_31_AWLOCK;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [2:0] m_axi_in_31_AWPROT;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [3:0] m_axi_in_31_AWQOS;
  (* RS_HS = "m_axi_in_31_AW.ready" *)input m_axi_in_31_AWREADY;
  (* RS_HS = "m_axi_in_31_AW.data" *)output [2:0] m_axi_in_31_AWSIZE;
  (* RS_HS = "m_axi_in_31_AW.valid" *)output m_axi_in_31_AWVALID;
  (* RS_HS = "m_axi_in_31_B.data" *)input [0:0] m_axi_in_31_BID;
  (* RS_HS = "m_axi_in_31_B.ready" *)output m_axi_in_31_BREADY;
  (* RS_HS = "m_axi_in_31_B.data" *)input [1:0] m_axi_in_31_BRESP;
  (* RS_HS = "m_axi_in_31_B.valid" *)input m_axi_in_31_BVALID;
  (* RS_HS = "m_axi_in_31_R.data" *)input [255:0] m_axi_in_31_RDATA;
  (* RS_HS = "m_axi_in_31_R.data" *)input [0:0] m_axi_in_31_RID;
  (* RS_HS = "m_axi_in_31_R.data" *)input m_axi_in_31_RLAST;
  (* RS_HS = "m_axi_in_31_R.ready" *)output m_axi_in_31_RREADY;
  (* RS_HS = "m_axi_in_31_R.data" *)input [1:0] m_axi_in_31_RRESP;
  (* RS_HS = "m_axi_in_31_R.valid" *)input m_axi_in_31_RVALID;
  (* RS_HS = "m_axi_in_31_W.data" *)output [255:0] m_axi_in_31_WDATA;
  (* RS_HS = "m_axi_in_31_W.data" *)output m_axi_in_31_WLAST;
  (* RS_HS = "m_axi_in_31_W.ready" *)input m_axi_in_31_WREADY;
  (* RS_HS = "m_axi_in_31_W.data" *)output [31:0] m_axi_in_31_WSTRB;
  (* RS_HS = "m_axi_in_31_W.valid" *)output m_axi_in_31_WVALID;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [63:0] m_axi_in_32_ARADDR;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [1:0] m_axi_in_32_ARBURST;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [3:0] m_axi_in_32_ARCACHE;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [0:0] m_axi_in_32_ARID;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [7:0] m_axi_in_32_ARLEN;
  (* RS_HS = "m_axi_in_32_AR.data" *)output m_axi_in_32_ARLOCK;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [2:0] m_axi_in_32_ARPROT;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [3:0] m_axi_in_32_ARQOS;
  (* RS_HS = "m_axi_in_32_AR.ready" *)input m_axi_in_32_ARREADY;
  (* RS_HS = "m_axi_in_32_AR.data" *)output [2:0] m_axi_in_32_ARSIZE;
  (* RS_HS = "m_axi_in_32_AR.valid" *)output m_axi_in_32_ARVALID;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [63:0] m_axi_in_32_AWADDR;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [1:0] m_axi_in_32_AWBURST;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [3:0] m_axi_in_32_AWCACHE;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [0:0] m_axi_in_32_AWID;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [7:0] m_axi_in_32_AWLEN;
  (* RS_HS = "m_axi_in_32_AW.data" *)output m_axi_in_32_AWLOCK;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [2:0] m_axi_in_32_AWPROT;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [3:0] m_axi_in_32_AWQOS;
  (* RS_HS = "m_axi_in_32_AW.ready" *)input m_axi_in_32_AWREADY;
  (* RS_HS = "m_axi_in_32_AW.data" *)output [2:0] m_axi_in_32_AWSIZE;
  (* RS_HS = "m_axi_in_32_AW.valid" *)output m_axi_in_32_AWVALID;
  (* RS_HS = "m_axi_in_32_B.data" *)input [0:0] m_axi_in_32_BID;
  (* RS_HS = "m_axi_in_32_B.ready" *)output m_axi_in_32_BREADY;
  (* RS_HS = "m_axi_in_32_B.data" *)input [1:0] m_axi_in_32_BRESP;
  (* RS_HS = "m_axi_in_32_B.valid" *)input m_axi_in_32_BVALID;
  (* RS_HS = "m_axi_in_32_R.data" *)input [255:0] m_axi_in_32_RDATA;
  (* RS_HS = "m_axi_in_32_R.data" *)input [0:0] m_axi_in_32_RID;
  (* RS_HS = "m_axi_in_32_R.data" *)input m_axi_in_32_RLAST;
  (* RS_HS = "m_axi_in_32_R.ready" *)output m_axi_in_32_RREADY;
  (* RS_HS = "m_axi_in_32_R.data" *)input [1:0] m_axi_in_32_RRESP;
  (* RS_HS = "m_axi_in_32_R.valid" *)input m_axi_in_32_RVALID;
  (* RS_HS = "m_axi_in_32_W.data" *)output [255:0] m_axi_in_32_WDATA;
  (* RS_HS = "m_axi_in_32_W.data" *)output m_axi_in_32_WLAST;
  (* RS_HS = "m_axi_in_32_W.ready" *)input m_axi_in_32_WREADY;
  (* RS_HS = "m_axi_in_32_W.data" *)output [31:0] m_axi_in_32_WSTRB;
  (* RS_HS = "m_axi_in_32_W.valid" *)output m_axi_in_32_WVALID;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [63:0] m_axi_in_33_ARADDR;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [1:0] m_axi_in_33_ARBURST;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [3:0] m_axi_in_33_ARCACHE;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [0:0] m_axi_in_33_ARID;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [7:0] m_axi_in_33_ARLEN;
  (* RS_HS = "m_axi_in_33_AR.data" *)output m_axi_in_33_ARLOCK;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [2:0] m_axi_in_33_ARPROT;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [3:0] m_axi_in_33_ARQOS;
  (* RS_HS = "m_axi_in_33_AR.ready" *)input m_axi_in_33_ARREADY;
  (* RS_HS = "m_axi_in_33_AR.data" *)output [2:0] m_axi_in_33_ARSIZE;
  (* RS_HS = "m_axi_in_33_AR.valid" *)output m_axi_in_33_ARVALID;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [63:0] m_axi_in_33_AWADDR;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [1:0] m_axi_in_33_AWBURST;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [3:0] m_axi_in_33_AWCACHE;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [0:0] m_axi_in_33_AWID;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [7:0] m_axi_in_33_AWLEN;
  (* RS_HS = "m_axi_in_33_AW.data" *)output m_axi_in_33_AWLOCK;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [2:0] m_axi_in_33_AWPROT;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [3:0] m_axi_in_33_AWQOS;
  (* RS_HS = "m_axi_in_33_AW.ready" *)input m_axi_in_33_AWREADY;
  (* RS_HS = "m_axi_in_33_AW.data" *)output [2:0] m_axi_in_33_AWSIZE;
  (* RS_HS = "m_axi_in_33_AW.valid" *)output m_axi_in_33_AWVALID;
  (* RS_HS = "m_axi_in_33_B.data" *)input [0:0] m_axi_in_33_BID;
  (* RS_HS = "m_axi_in_33_B.ready" *)output m_axi_in_33_BREADY;
  (* RS_HS = "m_axi_in_33_B.data" *)input [1:0] m_axi_in_33_BRESP;
  (* RS_HS = "m_axi_in_33_B.valid" *)input m_axi_in_33_BVALID;
  (* RS_HS = "m_axi_in_33_R.data" *)input [255:0] m_axi_in_33_RDATA;
  (* RS_HS = "m_axi_in_33_R.data" *)input [0:0] m_axi_in_33_RID;
  (* RS_HS = "m_axi_in_33_R.data" *)input m_axi_in_33_RLAST;
  (* RS_HS = "m_axi_in_33_R.ready" *)output m_axi_in_33_RREADY;
  (* RS_HS = "m_axi_in_33_R.data" *)input [1:0] m_axi_in_33_RRESP;
  (* RS_HS = "m_axi_in_33_R.valid" *)input m_axi_in_33_RVALID;
  (* RS_HS = "m_axi_in_33_W.data" *)output [255:0] m_axi_in_33_WDATA;
  (* RS_HS = "m_axi_in_33_W.data" *)output m_axi_in_33_WLAST;
  (* RS_HS = "m_axi_in_33_W.ready" *)input m_axi_in_33_WREADY;
  (* RS_HS = "m_axi_in_33_W.data" *)output [31:0] m_axi_in_33_WSTRB;
  (* RS_HS = "m_axi_in_33_W.valid" *)output m_axi_in_33_WVALID;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [63:0] m_axi_in_34_ARADDR;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [1:0] m_axi_in_34_ARBURST;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [3:0] m_axi_in_34_ARCACHE;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [0:0] m_axi_in_34_ARID;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [7:0] m_axi_in_34_ARLEN;
  (* RS_HS = "m_axi_in_34_AR.data" *)output m_axi_in_34_ARLOCK;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [2:0] m_axi_in_34_ARPROT;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [3:0] m_axi_in_34_ARQOS;
  (* RS_HS = "m_axi_in_34_AR.ready" *)input m_axi_in_34_ARREADY;
  (* RS_HS = "m_axi_in_34_AR.data" *)output [2:0] m_axi_in_34_ARSIZE;
  (* RS_HS = "m_axi_in_34_AR.valid" *)output m_axi_in_34_ARVALID;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [63:0] m_axi_in_34_AWADDR;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [1:0] m_axi_in_34_AWBURST;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [3:0] m_axi_in_34_AWCACHE;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [0:0] m_axi_in_34_AWID;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [7:0] m_axi_in_34_AWLEN;
  (* RS_HS = "m_axi_in_34_AW.data" *)output m_axi_in_34_AWLOCK;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [2:0] m_axi_in_34_AWPROT;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [3:0] m_axi_in_34_AWQOS;
  (* RS_HS = "m_axi_in_34_AW.ready" *)input m_axi_in_34_AWREADY;
  (* RS_HS = "m_axi_in_34_AW.data" *)output [2:0] m_axi_in_34_AWSIZE;
  (* RS_HS = "m_axi_in_34_AW.valid" *)output m_axi_in_34_AWVALID;
  (* RS_HS = "m_axi_in_34_B.data" *)input [0:0] m_axi_in_34_BID;
  (* RS_HS = "m_axi_in_34_B.ready" *)output m_axi_in_34_BREADY;
  (* RS_HS = "m_axi_in_34_B.data" *)input [1:0] m_axi_in_34_BRESP;
  (* RS_HS = "m_axi_in_34_B.valid" *)input m_axi_in_34_BVALID;
  (* RS_HS = "m_axi_in_34_R.data" *)input [255:0] m_axi_in_34_RDATA;
  (* RS_HS = "m_axi_in_34_R.data" *)input [0:0] m_axi_in_34_RID;
  (* RS_HS = "m_axi_in_34_R.data" *)input m_axi_in_34_RLAST;
  (* RS_HS = "m_axi_in_34_R.ready" *)output m_axi_in_34_RREADY;
  (* RS_HS = "m_axi_in_34_R.data" *)input [1:0] m_axi_in_34_RRESP;
  (* RS_HS = "m_axi_in_34_R.valid" *)input m_axi_in_34_RVALID;
  (* RS_HS = "m_axi_in_34_W.data" *)output [255:0] m_axi_in_34_WDATA;
  (* RS_HS = "m_axi_in_34_W.data" *)output m_axi_in_34_WLAST;
  (* RS_HS = "m_axi_in_34_W.ready" *)input m_axi_in_34_WREADY;
  (* RS_HS = "m_axi_in_34_W.data" *)output [31:0] m_axi_in_34_WSTRB;
  (* RS_HS = "m_axi_in_34_W.valid" *)output m_axi_in_34_WVALID;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [63:0] m_axi_in_35_ARADDR;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [1:0] m_axi_in_35_ARBURST;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [3:0] m_axi_in_35_ARCACHE;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [0:0] m_axi_in_35_ARID;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [7:0] m_axi_in_35_ARLEN;
  (* RS_HS = "m_axi_in_35_AR.data" *)output m_axi_in_35_ARLOCK;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [2:0] m_axi_in_35_ARPROT;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [3:0] m_axi_in_35_ARQOS;
  (* RS_HS = "m_axi_in_35_AR.ready" *)input m_axi_in_35_ARREADY;
  (* RS_HS = "m_axi_in_35_AR.data" *)output [2:0] m_axi_in_35_ARSIZE;
  (* RS_HS = "m_axi_in_35_AR.valid" *)output m_axi_in_35_ARVALID;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [63:0] m_axi_in_35_AWADDR;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [1:0] m_axi_in_35_AWBURST;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [3:0] m_axi_in_35_AWCACHE;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [0:0] m_axi_in_35_AWID;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [7:0] m_axi_in_35_AWLEN;
  (* RS_HS = "m_axi_in_35_AW.data" *)output m_axi_in_35_AWLOCK;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [2:0] m_axi_in_35_AWPROT;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [3:0] m_axi_in_35_AWQOS;
  (* RS_HS = "m_axi_in_35_AW.ready" *)input m_axi_in_35_AWREADY;
  (* RS_HS = "m_axi_in_35_AW.data" *)output [2:0] m_axi_in_35_AWSIZE;
  (* RS_HS = "m_axi_in_35_AW.valid" *)output m_axi_in_35_AWVALID;
  (* RS_HS = "m_axi_in_35_B.data" *)input [0:0] m_axi_in_35_BID;
  (* RS_HS = "m_axi_in_35_B.ready" *)output m_axi_in_35_BREADY;
  (* RS_HS = "m_axi_in_35_B.data" *)input [1:0] m_axi_in_35_BRESP;
  (* RS_HS = "m_axi_in_35_B.valid" *)input m_axi_in_35_BVALID;
  (* RS_HS = "m_axi_in_35_R.data" *)input [255:0] m_axi_in_35_RDATA;
  (* RS_HS = "m_axi_in_35_R.data" *)input [0:0] m_axi_in_35_RID;
  (* RS_HS = "m_axi_in_35_R.data" *)input m_axi_in_35_RLAST;
  (* RS_HS = "m_axi_in_35_R.ready" *)output m_axi_in_35_RREADY;
  (* RS_HS = "m_axi_in_35_R.data" *)input [1:0] m_axi_in_35_RRESP;
  (* RS_HS = "m_axi_in_35_R.valid" *)input m_axi_in_35_RVALID;
  (* RS_HS = "m_axi_in_35_W.data" *)output [255:0] m_axi_in_35_WDATA;
  (* RS_HS = "m_axi_in_35_W.data" *)output m_axi_in_35_WLAST;
  (* RS_HS = "m_axi_in_35_W.ready" *)input m_axi_in_35_WREADY;
  (* RS_HS = "m_axi_in_35_W.data" *)output [31:0] m_axi_in_35_WSTRB;
  (* RS_HS = "m_axi_in_35_W.valid" *)output m_axi_in_35_WVALID;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [63:0] m_axi_in_36_ARADDR;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [1:0] m_axi_in_36_ARBURST;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [3:0] m_axi_in_36_ARCACHE;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [0:0] m_axi_in_36_ARID;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [7:0] m_axi_in_36_ARLEN;
  (* RS_HS = "m_axi_in_36_AR.data" *)output m_axi_in_36_ARLOCK;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [2:0] m_axi_in_36_ARPROT;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [3:0] m_axi_in_36_ARQOS;
  (* RS_HS = "m_axi_in_36_AR.ready" *)input m_axi_in_36_ARREADY;
  (* RS_HS = "m_axi_in_36_AR.data" *)output [2:0] m_axi_in_36_ARSIZE;
  (* RS_HS = "m_axi_in_36_AR.valid" *)output m_axi_in_36_ARVALID;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [63:0] m_axi_in_36_AWADDR;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [1:0] m_axi_in_36_AWBURST;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [3:0] m_axi_in_36_AWCACHE;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [0:0] m_axi_in_36_AWID;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [7:0] m_axi_in_36_AWLEN;
  (* RS_HS = "m_axi_in_36_AW.data" *)output m_axi_in_36_AWLOCK;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [2:0] m_axi_in_36_AWPROT;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [3:0] m_axi_in_36_AWQOS;
  (* RS_HS = "m_axi_in_36_AW.ready" *)input m_axi_in_36_AWREADY;
  (* RS_HS = "m_axi_in_36_AW.data" *)output [2:0] m_axi_in_36_AWSIZE;
  (* RS_HS = "m_axi_in_36_AW.valid" *)output m_axi_in_36_AWVALID;
  (* RS_HS = "m_axi_in_36_B.data" *)input [0:0] m_axi_in_36_BID;
  (* RS_HS = "m_axi_in_36_B.ready" *)output m_axi_in_36_BREADY;
  (* RS_HS = "m_axi_in_36_B.data" *)input [1:0] m_axi_in_36_BRESP;
  (* RS_HS = "m_axi_in_36_B.valid" *)input m_axi_in_36_BVALID;
  (* RS_HS = "m_axi_in_36_R.data" *)input [255:0] m_axi_in_36_RDATA;
  (* RS_HS = "m_axi_in_36_R.data" *)input [0:0] m_axi_in_36_RID;
  (* RS_HS = "m_axi_in_36_R.data" *)input m_axi_in_36_RLAST;
  (* RS_HS = "m_axi_in_36_R.ready" *)output m_axi_in_36_RREADY;
  (* RS_HS = "m_axi_in_36_R.data" *)input [1:0] m_axi_in_36_RRESP;
  (* RS_HS = "m_axi_in_36_R.valid" *)input m_axi_in_36_RVALID;
  (* RS_HS = "m_axi_in_36_W.data" *)output [255:0] m_axi_in_36_WDATA;
  (* RS_HS = "m_axi_in_36_W.data" *)output m_axi_in_36_WLAST;
  (* RS_HS = "m_axi_in_36_W.ready" *)input m_axi_in_36_WREADY;
  (* RS_HS = "m_axi_in_36_W.data" *)output [31:0] m_axi_in_36_WSTRB;
  (* RS_HS = "m_axi_in_36_W.valid" *)output m_axi_in_36_WVALID;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [63:0] m_axi_in_37_ARADDR;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [1:0] m_axi_in_37_ARBURST;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [3:0] m_axi_in_37_ARCACHE;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [0:0] m_axi_in_37_ARID;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [7:0] m_axi_in_37_ARLEN;
  (* RS_HS = "m_axi_in_37_AR.data" *)output m_axi_in_37_ARLOCK;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [2:0] m_axi_in_37_ARPROT;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [3:0] m_axi_in_37_ARQOS;
  (* RS_HS = "m_axi_in_37_AR.ready" *)input m_axi_in_37_ARREADY;
  (* RS_HS = "m_axi_in_37_AR.data" *)output [2:0] m_axi_in_37_ARSIZE;
  (* RS_HS = "m_axi_in_37_AR.valid" *)output m_axi_in_37_ARVALID;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [63:0] m_axi_in_37_AWADDR;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [1:0] m_axi_in_37_AWBURST;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [3:0] m_axi_in_37_AWCACHE;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [0:0] m_axi_in_37_AWID;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [7:0] m_axi_in_37_AWLEN;
  (* RS_HS = "m_axi_in_37_AW.data" *)output m_axi_in_37_AWLOCK;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [2:0] m_axi_in_37_AWPROT;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [3:0] m_axi_in_37_AWQOS;
  (* RS_HS = "m_axi_in_37_AW.ready" *)input m_axi_in_37_AWREADY;
  (* RS_HS = "m_axi_in_37_AW.data" *)output [2:0] m_axi_in_37_AWSIZE;
  (* RS_HS = "m_axi_in_37_AW.valid" *)output m_axi_in_37_AWVALID;
  (* RS_HS = "m_axi_in_37_B.data" *)input [0:0] m_axi_in_37_BID;
  (* RS_HS = "m_axi_in_37_B.ready" *)output m_axi_in_37_BREADY;
  (* RS_HS = "m_axi_in_37_B.data" *)input [1:0] m_axi_in_37_BRESP;
  (* RS_HS = "m_axi_in_37_B.valid" *)input m_axi_in_37_BVALID;
  (* RS_HS = "m_axi_in_37_R.data" *)input [255:0] m_axi_in_37_RDATA;
  (* RS_HS = "m_axi_in_37_R.data" *)input [0:0] m_axi_in_37_RID;
  (* RS_HS = "m_axi_in_37_R.data" *)input m_axi_in_37_RLAST;
  (* RS_HS = "m_axi_in_37_R.ready" *)output m_axi_in_37_RREADY;
  (* RS_HS = "m_axi_in_37_R.data" *)input [1:0] m_axi_in_37_RRESP;
  (* RS_HS = "m_axi_in_37_R.valid" *)input m_axi_in_37_RVALID;
  (* RS_HS = "m_axi_in_37_W.data" *)output [255:0] m_axi_in_37_WDATA;
  (* RS_HS = "m_axi_in_37_W.data" *)output m_axi_in_37_WLAST;
  (* RS_HS = "m_axi_in_37_W.ready" *)input m_axi_in_37_WREADY;
  (* RS_HS = "m_axi_in_37_W.data" *)output [31:0] m_axi_in_37_WSTRB;
  (* RS_HS = "m_axi_in_37_W.valid" *)output m_axi_in_37_WVALID;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [63:0] m_axi_in_38_ARADDR;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [1:0] m_axi_in_38_ARBURST;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [3:0] m_axi_in_38_ARCACHE;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [0:0] m_axi_in_38_ARID;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [7:0] m_axi_in_38_ARLEN;
  (* RS_HS = "m_axi_in_38_AR.data" *)output m_axi_in_38_ARLOCK;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [2:0] m_axi_in_38_ARPROT;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [3:0] m_axi_in_38_ARQOS;
  (* RS_HS = "m_axi_in_38_AR.ready" *)input m_axi_in_38_ARREADY;
  (* RS_HS = "m_axi_in_38_AR.data" *)output [2:0] m_axi_in_38_ARSIZE;
  (* RS_HS = "m_axi_in_38_AR.valid" *)output m_axi_in_38_ARVALID;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [63:0] m_axi_in_38_AWADDR;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [1:0] m_axi_in_38_AWBURST;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [3:0] m_axi_in_38_AWCACHE;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [0:0] m_axi_in_38_AWID;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [7:0] m_axi_in_38_AWLEN;
  (* RS_HS = "m_axi_in_38_AW.data" *)output m_axi_in_38_AWLOCK;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [2:0] m_axi_in_38_AWPROT;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [3:0] m_axi_in_38_AWQOS;
  (* RS_HS = "m_axi_in_38_AW.ready" *)input m_axi_in_38_AWREADY;
  (* RS_HS = "m_axi_in_38_AW.data" *)output [2:0] m_axi_in_38_AWSIZE;
  (* RS_HS = "m_axi_in_38_AW.valid" *)output m_axi_in_38_AWVALID;
  (* RS_HS = "m_axi_in_38_B.data" *)input [0:0] m_axi_in_38_BID;
  (* RS_HS = "m_axi_in_38_B.ready" *)output m_axi_in_38_BREADY;
  (* RS_HS = "m_axi_in_38_B.data" *)input [1:0] m_axi_in_38_BRESP;
  (* RS_HS = "m_axi_in_38_B.valid" *)input m_axi_in_38_BVALID;
  (* RS_HS = "m_axi_in_38_R.data" *)input [255:0] m_axi_in_38_RDATA;
  (* RS_HS = "m_axi_in_38_R.data" *)input [0:0] m_axi_in_38_RID;
  (* RS_HS = "m_axi_in_38_R.data" *)input m_axi_in_38_RLAST;
  (* RS_HS = "m_axi_in_38_R.ready" *)output m_axi_in_38_RREADY;
  (* RS_HS = "m_axi_in_38_R.data" *)input [1:0] m_axi_in_38_RRESP;
  (* RS_HS = "m_axi_in_38_R.valid" *)input m_axi_in_38_RVALID;
  (* RS_HS = "m_axi_in_38_W.data" *)output [255:0] m_axi_in_38_WDATA;
  (* RS_HS = "m_axi_in_38_W.data" *)output m_axi_in_38_WLAST;
  (* RS_HS = "m_axi_in_38_W.ready" *)input m_axi_in_38_WREADY;
  (* RS_HS = "m_axi_in_38_W.data" *)output [31:0] m_axi_in_38_WSTRB;
  (* RS_HS = "m_axi_in_38_W.valid" *)output m_axi_in_38_WVALID;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [63:0] m_axi_in_39_ARADDR;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [1:0] m_axi_in_39_ARBURST;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [3:0] m_axi_in_39_ARCACHE;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [0:0] m_axi_in_39_ARID;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [7:0] m_axi_in_39_ARLEN;
  (* RS_HS = "m_axi_in_39_AR.data" *)output m_axi_in_39_ARLOCK;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [2:0] m_axi_in_39_ARPROT;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [3:0] m_axi_in_39_ARQOS;
  (* RS_HS = "m_axi_in_39_AR.ready" *)input m_axi_in_39_ARREADY;
  (* RS_HS = "m_axi_in_39_AR.data" *)output [2:0] m_axi_in_39_ARSIZE;
  (* RS_HS = "m_axi_in_39_AR.valid" *)output m_axi_in_39_ARVALID;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [63:0] m_axi_in_39_AWADDR;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [1:0] m_axi_in_39_AWBURST;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [3:0] m_axi_in_39_AWCACHE;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [0:0] m_axi_in_39_AWID;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [7:0] m_axi_in_39_AWLEN;
  (* RS_HS = "m_axi_in_39_AW.data" *)output m_axi_in_39_AWLOCK;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [2:0] m_axi_in_39_AWPROT;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [3:0] m_axi_in_39_AWQOS;
  (* RS_HS = "m_axi_in_39_AW.ready" *)input m_axi_in_39_AWREADY;
  (* RS_HS = "m_axi_in_39_AW.data" *)output [2:0] m_axi_in_39_AWSIZE;
  (* RS_HS = "m_axi_in_39_AW.valid" *)output m_axi_in_39_AWVALID;
  (* RS_HS = "m_axi_in_39_B.data" *)input [0:0] m_axi_in_39_BID;
  (* RS_HS = "m_axi_in_39_B.ready" *)output m_axi_in_39_BREADY;
  (* RS_HS = "m_axi_in_39_B.data" *)input [1:0] m_axi_in_39_BRESP;
  (* RS_HS = "m_axi_in_39_B.valid" *)input m_axi_in_39_BVALID;
  (* RS_HS = "m_axi_in_39_R.data" *)input [255:0] m_axi_in_39_RDATA;
  (* RS_HS = "m_axi_in_39_R.data" *)input [0:0] m_axi_in_39_RID;
  (* RS_HS = "m_axi_in_39_R.data" *)input m_axi_in_39_RLAST;
  (* RS_HS = "m_axi_in_39_R.ready" *)output m_axi_in_39_RREADY;
  (* RS_HS = "m_axi_in_39_R.data" *)input [1:0] m_axi_in_39_RRESP;
  (* RS_HS = "m_axi_in_39_R.valid" *)input m_axi_in_39_RVALID;
  (* RS_HS = "m_axi_in_39_W.data" *)output [255:0] m_axi_in_39_WDATA;
  (* RS_HS = "m_axi_in_39_W.data" *)output m_axi_in_39_WLAST;
  (* RS_HS = "m_axi_in_39_W.ready" *)input m_axi_in_39_WREADY;
  (* RS_HS = "m_axi_in_39_W.data" *)output [31:0] m_axi_in_39_WSTRB;
  (* RS_HS = "m_axi_in_39_W.valid" *)output m_axi_in_39_WVALID;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [63:0] m_axi_in_4_ARADDR;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [1:0] m_axi_in_4_ARBURST;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [3:0] m_axi_in_4_ARCACHE;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [0:0] m_axi_in_4_ARID;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [7:0] m_axi_in_4_ARLEN;
  (* RS_HS = "m_axi_in_4_AR.data" *)output m_axi_in_4_ARLOCK;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [2:0] m_axi_in_4_ARPROT;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [3:0] m_axi_in_4_ARQOS;
  (* RS_HS = "m_axi_in_4_AR.ready" *)input m_axi_in_4_ARREADY;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [2:0] m_axi_in_4_ARSIZE;
  (* RS_HS = "m_axi_in_4_AR.valid" *)output m_axi_in_4_ARVALID;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [63:0] m_axi_in_4_AWADDR;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [1:0] m_axi_in_4_AWBURST;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [3:0] m_axi_in_4_AWCACHE;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [0:0] m_axi_in_4_AWID;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [7:0] m_axi_in_4_AWLEN;
  (* RS_HS = "m_axi_in_4_AW.data" *)output m_axi_in_4_AWLOCK;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [2:0] m_axi_in_4_AWPROT;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [3:0] m_axi_in_4_AWQOS;
  (* RS_HS = "m_axi_in_4_AW.ready" *)input m_axi_in_4_AWREADY;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [2:0] m_axi_in_4_AWSIZE;
  (* RS_HS = "m_axi_in_4_AW.valid" *)output m_axi_in_4_AWVALID;
  (* RS_HS = "m_axi_in_4_B.data" *)input [0:0] m_axi_in_4_BID;
  (* RS_HS = "m_axi_in_4_B.ready" *)output m_axi_in_4_BREADY;
  (* RS_HS = "m_axi_in_4_B.data" *)input [1:0] m_axi_in_4_BRESP;
  (* RS_HS = "m_axi_in_4_B.valid" *)input m_axi_in_4_BVALID;
  (* RS_HS = "m_axi_in_4_R.data" *)input [255:0] m_axi_in_4_RDATA;
  (* RS_HS = "m_axi_in_4_R.data" *)input [0:0] m_axi_in_4_RID;
  (* RS_HS = "m_axi_in_4_R.data" *)input m_axi_in_4_RLAST;
  (* RS_HS = "m_axi_in_4_R.ready" *)output m_axi_in_4_RREADY;
  (* RS_HS = "m_axi_in_4_R.data" *)input [1:0] m_axi_in_4_RRESP;
  (* RS_HS = "m_axi_in_4_R.valid" *)input m_axi_in_4_RVALID;
  (* RS_HS = "m_axi_in_4_W.data" *)output [255:0] m_axi_in_4_WDATA;
  (* RS_HS = "m_axi_in_4_W.data" *)output m_axi_in_4_WLAST;
  (* RS_HS = "m_axi_in_4_W.ready" *)input m_axi_in_4_WREADY;
  (* RS_HS = "m_axi_in_4_W.data" *)output [31:0] m_axi_in_4_WSTRB;
  (* RS_HS = "m_axi_in_4_W.valid" *)output m_axi_in_4_WVALID;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [63:0] m_axi_in_40_ARADDR;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [1:0] m_axi_in_40_ARBURST;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [3:0] m_axi_in_40_ARCACHE;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [0:0] m_axi_in_40_ARID;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [7:0] m_axi_in_40_ARLEN;
  (* RS_HS = "m_axi_in_40_AR.data" *)output m_axi_in_40_ARLOCK;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [2:0] m_axi_in_40_ARPROT;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [3:0] m_axi_in_40_ARQOS;
  (* RS_HS = "m_axi_in_40_AR.ready" *)input m_axi_in_40_ARREADY;
  (* RS_HS = "m_axi_in_40_AR.data" *)output [2:0] m_axi_in_40_ARSIZE;
  (* RS_HS = "m_axi_in_40_AR.valid" *)output m_axi_in_40_ARVALID;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [63:0] m_axi_in_40_AWADDR;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [1:0] m_axi_in_40_AWBURST;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [3:0] m_axi_in_40_AWCACHE;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [0:0] m_axi_in_40_AWID;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [7:0] m_axi_in_40_AWLEN;
  (* RS_HS = "m_axi_in_40_AW.data" *)output m_axi_in_40_AWLOCK;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [2:0] m_axi_in_40_AWPROT;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [3:0] m_axi_in_40_AWQOS;
  (* RS_HS = "m_axi_in_40_AW.ready" *)input m_axi_in_40_AWREADY;
  (* RS_HS = "m_axi_in_40_AW.data" *)output [2:0] m_axi_in_40_AWSIZE;
  (* RS_HS = "m_axi_in_40_AW.valid" *)output m_axi_in_40_AWVALID;
  (* RS_HS = "m_axi_in_40_B.data" *)input [0:0] m_axi_in_40_BID;
  (* RS_HS = "m_axi_in_40_B.ready" *)output m_axi_in_40_BREADY;
  (* RS_HS = "m_axi_in_40_B.data" *)input [1:0] m_axi_in_40_BRESP;
  (* RS_HS = "m_axi_in_40_B.valid" *)input m_axi_in_40_BVALID;
  (* RS_HS = "m_axi_in_40_R.data" *)input [255:0] m_axi_in_40_RDATA;
  (* RS_HS = "m_axi_in_40_R.data" *)input [0:0] m_axi_in_40_RID;
  (* RS_HS = "m_axi_in_40_R.data" *)input m_axi_in_40_RLAST;
  (* RS_HS = "m_axi_in_40_R.ready" *)output m_axi_in_40_RREADY;
  (* RS_HS = "m_axi_in_40_R.data" *)input [1:0] m_axi_in_40_RRESP;
  (* RS_HS = "m_axi_in_40_R.valid" *)input m_axi_in_40_RVALID;
  (* RS_HS = "m_axi_in_40_W.data" *)output [255:0] m_axi_in_40_WDATA;
  (* RS_HS = "m_axi_in_40_W.data" *)output m_axi_in_40_WLAST;
  (* RS_HS = "m_axi_in_40_W.ready" *)input m_axi_in_40_WREADY;
  (* RS_HS = "m_axi_in_40_W.data" *)output [31:0] m_axi_in_40_WSTRB;
  (* RS_HS = "m_axi_in_40_W.valid" *)output m_axi_in_40_WVALID;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [63:0] m_axi_in_41_ARADDR;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [1:0] m_axi_in_41_ARBURST;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [3:0] m_axi_in_41_ARCACHE;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [0:0] m_axi_in_41_ARID;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [7:0] m_axi_in_41_ARLEN;
  (* RS_HS = "m_axi_in_41_AR.data" *)output m_axi_in_41_ARLOCK;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [2:0] m_axi_in_41_ARPROT;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [3:0] m_axi_in_41_ARQOS;
  (* RS_HS = "m_axi_in_41_AR.ready" *)input m_axi_in_41_ARREADY;
  (* RS_HS = "m_axi_in_41_AR.data" *)output [2:0] m_axi_in_41_ARSIZE;
  (* RS_HS = "m_axi_in_41_AR.valid" *)output m_axi_in_41_ARVALID;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [63:0] m_axi_in_41_AWADDR;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [1:0] m_axi_in_41_AWBURST;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [3:0] m_axi_in_41_AWCACHE;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [0:0] m_axi_in_41_AWID;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [7:0] m_axi_in_41_AWLEN;
  (* RS_HS = "m_axi_in_41_AW.data" *)output m_axi_in_41_AWLOCK;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [2:0] m_axi_in_41_AWPROT;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [3:0] m_axi_in_41_AWQOS;
  (* RS_HS = "m_axi_in_41_AW.ready" *)input m_axi_in_41_AWREADY;
  (* RS_HS = "m_axi_in_41_AW.data" *)output [2:0] m_axi_in_41_AWSIZE;
  (* RS_HS = "m_axi_in_41_AW.valid" *)output m_axi_in_41_AWVALID;
  (* RS_HS = "m_axi_in_41_B.data" *)input [0:0] m_axi_in_41_BID;
  (* RS_HS = "m_axi_in_41_B.ready" *)output m_axi_in_41_BREADY;
  (* RS_HS = "m_axi_in_41_B.data" *)input [1:0] m_axi_in_41_BRESP;
  (* RS_HS = "m_axi_in_41_B.valid" *)input m_axi_in_41_BVALID;
  (* RS_HS = "m_axi_in_41_R.data" *)input [255:0] m_axi_in_41_RDATA;
  (* RS_HS = "m_axi_in_41_R.data" *)input [0:0] m_axi_in_41_RID;
  (* RS_HS = "m_axi_in_41_R.data" *)input m_axi_in_41_RLAST;
  (* RS_HS = "m_axi_in_41_R.ready" *)output m_axi_in_41_RREADY;
  (* RS_HS = "m_axi_in_41_R.data" *)input [1:0] m_axi_in_41_RRESP;
  (* RS_HS = "m_axi_in_41_R.valid" *)input m_axi_in_41_RVALID;
  (* RS_HS = "m_axi_in_41_W.data" *)output [255:0] m_axi_in_41_WDATA;
  (* RS_HS = "m_axi_in_41_W.data" *)output m_axi_in_41_WLAST;
  (* RS_HS = "m_axi_in_41_W.ready" *)input m_axi_in_41_WREADY;
  (* RS_HS = "m_axi_in_41_W.data" *)output [31:0] m_axi_in_41_WSTRB;
  (* RS_HS = "m_axi_in_41_W.valid" *)output m_axi_in_41_WVALID;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [63:0] m_axi_in_42_ARADDR;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [1:0] m_axi_in_42_ARBURST;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [3:0] m_axi_in_42_ARCACHE;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [0:0] m_axi_in_42_ARID;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [7:0] m_axi_in_42_ARLEN;
  (* RS_HS = "m_axi_in_42_AR.data" *)output m_axi_in_42_ARLOCK;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [2:0] m_axi_in_42_ARPROT;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [3:0] m_axi_in_42_ARQOS;
  (* RS_HS = "m_axi_in_42_AR.ready" *)input m_axi_in_42_ARREADY;
  (* RS_HS = "m_axi_in_42_AR.data" *)output [2:0] m_axi_in_42_ARSIZE;
  (* RS_HS = "m_axi_in_42_AR.valid" *)output m_axi_in_42_ARVALID;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [63:0] m_axi_in_42_AWADDR;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [1:0] m_axi_in_42_AWBURST;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [3:0] m_axi_in_42_AWCACHE;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [0:0] m_axi_in_42_AWID;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [7:0] m_axi_in_42_AWLEN;
  (* RS_HS = "m_axi_in_42_AW.data" *)output m_axi_in_42_AWLOCK;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [2:0] m_axi_in_42_AWPROT;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [3:0] m_axi_in_42_AWQOS;
  (* RS_HS = "m_axi_in_42_AW.ready" *)input m_axi_in_42_AWREADY;
  (* RS_HS = "m_axi_in_42_AW.data" *)output [2:0] m_axi_in_42_AWSIZE;
  (* RS_HS = "m_axi_in_42_AW.valid" *)output m_axi_in_42_AWVALID;
  (* RS_HS = "m_axi_in_42_B.data" *)input [0:0] m_axi_in_42_BID;
  (* RS_HS = "m_axi_in_42_B.ready" *)output m_axi_in_42_BREADY;
  (* RS_HS = "m_axi_in_42_B.data" *)input [1:0] m_axi_in_42_BRESP;
  (* RS_HS = "m_axi_in_42_B.valid" *)input m_axi_in_42_BVALID;
  (* RS_HS = "m_axi_in_42_R.data" *)input [255:0] m_axi_in_42_RDATA;
  (* RS_HS = "m_axi_in_42_R.data" *)input [0:0] m_axi_in_42_RID;
  (* RS_HS = "m_axi_in_42_R.data" *)input m_axi_in_42_RLAST;
  (* RS_HS = "m_axi_in_42_R.ready" *)output m_axi_in_42_RREADY;
  (* RS_HS = "m_axi_in_42_R.data" *)input [1:0] m_axi_in_42_RRESP;
  (* RS_HS = "m_axi_in_42_R.valid" *)input m_axi_in_42_RVALID;
  (* RS_HS = "m_axi_in_42_W.data" *)output [255:0] m_axi_in_42_WDATA;
  (* RS_HS = "m_axi_in_42_W.data" *)output m_axi_in_42_WLAST;
  (* RS_HS = "m_axi_in_42_W.ready" *)input m_axi_in_42_WREADY;
  (* RS_HS = "m_axi_in_42_W.data" *)output [31:0] m_axi_in_42_WSTRB;
  (* RS_HS = "m_axi_in_42_W.valid" *)output m_axi_in_42_WVALID;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [63:0] m_axi_in_43_ARADDR;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [1:0] m_axi_in_43_ARBURST;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [3:0] m_axi_in_43_ARCACHE;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [0:0] m_axi_in_43_ARID;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [7:0] m_axi_in_43_ARLEN;
  (* RS_HS = "m_axi_in_43_AR.data" *)output m_axi_in_43_ARLOCK;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [2:0] m_axi_in_43_ARPROT;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [3:0] m_axi_in_43_ARQOS;
  (* RS_HS = "m_axi_in_43_AR.ready" *)input m_axi_in_43_ARREADY;
  (* RS_HS = "m_axi_in_43_AR.data" *)output [2:0] m_axi_in_43_ARSIZE;
  (* RS_HS = "m_axi_in_43_AR.valid" *)output m_axi_in_43_ARVALID;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [63:0] m_axi_in_43_AWADDR;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [1:0] m_axi_in_43_AWBURST;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [3:0] m_axi_in_43_AWCACHE;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [0:0] m_axi_in_43_AWID;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [7:0] m_axi_in_43_AWLEN;
  (* RS_HS = "m_axi_in_43_AW.data" *)output m_axi_in_43_AWLOCK;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [2:0] m_axi_in_43_AWPROT;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [3:0] m_axi_in_43_AWQOS;
  (* RS_HS = "m_axi_in_43_AW.ready" *)input m_axi_in_43_AWREADY;
  (* RS_HS = "m_axi_in_43_AW.data" *)output [2:0] m_axi_in_43_AWSIZE;
  (* RS_HS = "m_axi_in_43_AW.valid" *)output m_axi_in_43_AWVALID;
  (* RS_HS = "m_axi_in_43_B.data" *)input [0:0] m_axi_in_43_BID;
  (* RS_HS = "m_axi_in_43_B.ready" *)output m_axi_in_43_BREADY;
  (* RS_HS = "m_axi_in_43_B.data" *)input [1:0] m_axi_in_43_BRESP;
  (* RS_HS = "m_axi_in_43_B.valid" *)input m_axi_in_43_BVALID;
  (* RS_HS = "m_axi_in_43_R.data" *)input [255:0] m_axi_in_43_RDATA;
  (* RS_HS = "m_axi_in_43_R.data" *)input [0:0] m_axi_in_43_RID;
  (* RS_HS = "m_axi_in_43_R.data" *)input m_axi_in_43_RLAST;
  (* RS_HS = "m_axi_in_43_R.ready" *)output m_axi_in_43_RREADY;
  (* RS_HS = "m_axi_in_43_R.data" *)input [1:0] m_axi_in_43_RRESP;
  (* RS_HS = "m_axi_in_43_R.valid" *)input m_axi_in_43_RVALID;
  (* RS_HS = "m_axi_in_43_W.data" *)output [255:0] m_axi_in_43_WDATA;
  (* RS_HS = "m_axi_in_43_W.data" *)output m_axi_in_43_WLAST;
  (* RS_HS = "m_axi_in_43_W.ready" *)input m_axi_in_43_WREADY;
  (* RS_HS = "m_axi_in_43_W.data" *)output [31:0] m_axi_in_43_WSTRB;
  (* RS_HS = "m_axi_in_43_W.valid" *)output m_axi_in_43_WVALID;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [63:0] m_axi_in_44_ARADDR;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [1:0] m_axi_in_44_ARBURST;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [3:0] m_axi_in_44_ARCACHE;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [0:0] m_axi_in_44_ARID;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [7:0] m_axi_in_44_ARLEN;
  (* RS_HS = "m_axi_in_44_AR.data" *)output m_axi_in_44_ARLOCK;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [2:0] m_axi_in_44_ARPROT;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [3:0] m_axi_in_44_ARQOS;
  (* RS_HS = "m_axi_in_44_AR.ready" *)input m_axi_in_44_ARREADY;
  (* RS_HS = "m_axi_in_44_AR.data" *)output [2:0] m_axi_in_44_ARSIZE;
  (* RS_HS = "m_axi_in_44_AR.valid" *)output m_axi_in_44_ARVALID;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [63:0] m_axi_in_44_AWADDR;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [1:0] m_axi_in_44_AWBURST;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [3:0] m_axi_in_44_AWCACHE;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [0:0] m_axi_in_44_AWID;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [7:0] m_axi_in_44_AWLEN;
  (* RS_HS = "m_axi_in_44_AW.data" *)output m_axi_in_44_AWLOCK;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [2:0] m_axi_in_44_AWPROT;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [3:0] m_axi_in_44_AWQOS;
  (* RS_HS = "m_axi_in_44_AW.ready" *)input m_axi_in_44_AWREADY;
  (* RS_HS = "m_axi_in_44_AW.data" *)output [2:0] m_axi_in_44_AWSIZE;
  (* RS_HS = "m_axi_in_44_AW.valid" *)output m_axi_in_44_AWVALID;
  (* RS_HS = "m_axi_in_44_B.data" *)input [0:0] m_axi_in_44_BID;
  (* RS_HS = "m_axi_in_44_B.ready" *)output m_axi_in_44_BREADY;
  (* RS_HS = "m_axi_in_44_B.data" *)input [1:0] m_axi_in_44_BRESP;
  (* RS_HS = "m_axi_in_44_B.valid" *)input m_axi_in_44_BVALID;
  (* RS_HS = "m_axi_in_44_R.data" *)input [255:0] m_axi_in_44_RDATA;
  (* RS_HS = "m_axi_in_44_R.data" *)input [0:0] m_axi_in_44_RID;
  (* RS_HS = "m_axi_in_44_R.data" *)input m_axi_in_44_RLAST;
  (* RS_HS = "m_axi_in_44_R.ready" *)output m_axi_in_44_RREADY;
  (* RS_HS = "m_axi_in_44_R.data" *)input [1:0] m_axi_in_44_RRESP;
  (* RS_HS = "m_axi_in_44_R.valid" *)input m_axi_in_44_RVALID;
  (* RS_HS = "m_axi_in_44_W.data" *)output [255:0] m_axi_in_44_WDATA;
  (* RS_HS = "m_axi_in_44_W.data" *)output m_axi_in_44_WLAST;
  (* RS_HS = "m_axi_in_44_W.ready" *)input m_axi_in_44_WREADY;
  (* RS_HS = "m_axi_in_44_W.data" *)output [31:0] m_axi_in_44_WSTRB;
  (* RS_HS = "m_axi_in_44_W.valid" *)output m_axi_in_44_WVALID;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [63:0] m_axi_in_45_ARADDR;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [1:0] m_axi_in_45_ARBURST;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [3:0] m_axi_in_45_ARCACHE;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [0:0] m_axi_in_45_ARID;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [7:0] m_axi_in_45_ARLEN;
  (* RS_HS = "m_axi_in_45_AR.data" *)output m_axi_in_45_ARLOCK;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [2:0] m_axi_in_45_ARPROT;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [3:0] m_axi_in_45_ARQOS;
  (* RS_HS = "m_axi_in_45_AR.ready" *)input m_axi_in_45_ARREADY;
  (* RS_HS = "m_axi_in_45_AR.data" *)output [2:0] m_axi_in_45_ARSIZE;
  (* RS_HS = "m_axi_in_45_AR.valid" *)output m_axi_in_45_ARVALID;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [63:0] m_axi_in_45_AWADDR;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [1:0] m_axi_in_45_AWBURST;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [3:0] m_axi_in_45_AWCACHE;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [0:0] m_axi_in_45_AWID;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [7:0] m_axi_in_45_AWLEN;
  (* RS_HS = "m_axi_in_45_AW.data" *)output m_axi_in_45_AWLOCK;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [2:0] m_axi_in_45_AWPROT;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [3:0] m_axi_in_45_AWQOS;
  (* RS_HS = "m_axi_in_45_AW.ready" *)input m_axi_in_45_AWREADY;
  (* RS_HS = "m_axi_in_45_AW.data" *)output [2:0] m_axi_in_45_AWSIZE;
  (* RS_HS = "m_axi_in_45_AW.valid" *)output m_axi_in_45_AWVALID;
  (* RS_HS = "m_axi_in_45_B.data" *)input [0:0] m_axi_in_45_BID;
  (* RS_HS = "m_axi_in_45_B.ready" *)output m_axi_in_45_BREADY;
  (* RS_HS = "m_axi_in_45_B.data" *)input [1:0] m_axi_in_45_BRESP;
  (* RS_HS = "m_axi_in_45_B.valid" *)input m_axi_in_45_BVALID;
  (* RS_HS = "m_axi_in_45_R.data" *)input [255:0] m_axi_in_45_RDATA;
  (* RS_HS = "m_axi_in_45_R.data" *)input [0:0] m_axi_in_45_RID;
  (* RS_HS = "m_axi_in_45_R.data" *)input m_axi_in_45_RLAST;
  (* RS_HS = "m_axi_in_45_R.ready" *)output m_axi_in_45_RREADY;
  (* RS_HS = "m_axi_in_45_R.data" *)input [1:0] m_axi_in_45_RRESP;
  (* RS_HS = "m_axi_in_45_R.valid" *)input m_axi_in_45_RVALID;
  (* RS_HS = "m_axi_in_45_W.data" *)output [255:0] m_axi_in_45_WDATA;
  (* RS_HS = "m_axi_in_45_W.data" *)output m_axi_in_45_WLAST;
  (* RS_HS = "m_axi_in_45_W.ready" *)input m_axi_in_45_WREADY;
  (* RS_HS = "m_axi_in_45_W.data" *)output [31:0] m_axi_in_45_WSTRB;
  (* RS_HS = "m_axi_in_45_W.valid" *)output m_axi_in_45_WVALID;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [63:0] m_axi_in_46_ARADDR;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [1:0] m_axi_in_46_ARBURST;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [3:0] m_axi_in_46_ARCACHE;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [0:0] m_axi_in_46_ARID;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [7:0] m_axi_in_46_ARLEN;
  (* RS_HS = "m_axi_in_46_AR.data" *)output m_axi_in_46_ARLOCK;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [2:0] m_axi_in_46_ARPROT;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [3:0] m_axi_in_46_ARQOS;
  (* RS_HS = "m_axi_in_46_AR.ready" *)input m_axi_in_46_ARREADY;
  (* RS_HS = "m_axi_in_46_AR.data" *)output [2:0] m_axi_in_46_ARSIZE;
  (* RS_HS = "m_axi_in_46_AR.valid" *)output m_axi_in_46_ARVALID;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [63:0] m_axi_in_46_AWADDR;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [1:0] m_axi_in_46_AWBURST;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [3:0] m_axi_in_46_AWCACHE;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [0:0] m_axi_in_46_AWID;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [7:0] m_axi_in_46_AWLEN;
  (* RS_HS = "m_axi_in_46_AW.data" *)output m_axi_in_46_AWLOCK;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [2:0] m_axi_in_46_AWPROT;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [3:0] m_axi_in_46_AWQOS;
  (* RS_HS = "m_axi_in_46_AW.ready" *)input m_axi_in_46_AWREADY;
  (* RS_HS = "m_axi_in_46_AW.data" *)output [2:0] m_axi_in_46_AWSIZE;
  (* RS_HS = "m_axi_in_46_AW.valid" *)output m_axi_in_46_AWVALID;
  (* RS_HS = "m_axi_in_46_B.data" *)input [0:0] m_axi_in_46_BID;
  (* RS_HS = "m_axi_in_46_B.ready" *)output m_axi_in_46_BREADY;
  (* RS_HS = "m_axi_in_46_B.data" *)input [1:0] m_axi_in_46_BRESP;
  (* RS_HS = "m_axi_in_46_B.valid" *)input m_axi_in_46_BVALID;
  (* RS_HS = "m_axi_in_46_R.data" *)input [255:0] m_axi_in_46_RDATA;
  (* RS_HS = "m_axi_in_46_R.data" *)input [0:0] m_axi_in_46_RID;
  (* RS_HS = "m_axi_in_46_R.data" *)input m_axi_in_46_RLAST;
  (* RS_HS = "m_axi_in_46_R.ready" *)output m_axi_in_46_RREADY;
  (* RS_HS = "m_axi_in_46_R.data" *)input [1:0] m_axi_in_46_RRESP;
  (* RS_HS = "m_axi_in_46_R.valid" *)input m_axi_in_46_RVALID;
  (* RS_HS = "m_axi_in_46_W.data" *)output [255:0] m_axi_in_46_WDATA;
  (* RS_HS = "m_axi_in_46_W.data" *)output m_axi_in_46_WLAST;
  (* RS_HS = "m_axi_in_46_W.ready" *)input m_axi_in_46_WREADY;
  (* RS_HS = "m_axi_in_46_W.data" *)output [31:0] m_axi_in_46_WSTRB;
  (* RS_HS = "m_axi_in_46_W.valid" *)output m_axi_in_46_WVALID;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [63:0] m_axi_in_47_ARADDR;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [1:0] m_axi_in_47_ARBURST;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [3:0] m_axi_in_47_ARCACHE;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [0:0] m_axi_in_47_ARID;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [7:0] m_axi_in_47_ARLEN;
  (* RS_HS = "m_axi_in_47_AR.data" *)output m_axi_in_47_ARLOCK;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [2:0] m_axi_in_47_ARPROT;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [3:0] m_axi_in_47_ARQOS;
  (* RS_HS = "m_axi_in_47_AR.ready" *)input m_axi_in_47_ARREADY;
  (* RS_HS = "m_axi_in_47_AR.data" *)output [2:0] m_axi_in_47_ARSIZE;
  (* RS_HS = "m_axi_in_47_AR.valid" *)output m_axi_in_47_ARVALID;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [63:0] m_axi_in_47_AWADDR;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [1:0] m_axi_in_47_AWBURST;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [3:0] m_axi_in_47_AWCACHE;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [0:0] m_axi_in_47_AWID;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [7:0] m_axi_in_47_AWLEN;
  (* RS_HS = "m_axi_in_47_AW.data" *)output m_axi_in_47_AWLOCK;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [2:0] m_axi_in_47_AWPROT;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [3:0] m_axi_in_47_AWQOS;
  (* RS_HS = "m_axi_in_47_AW.ready" *)input m_axi_in_47_AWREADY;
  (* RS_HS = "m_axi_in_47_AW.data" *)output [2:0] m_axi_in_47_AWSIZE;
  (* RS_HS = "m_axi_in_47_AW.valid" *)output m_axi_in_47_AWVALID;
  (* RS_HS = "m_axi_in_47_B.data" *)input [0:0] m_axi_in_47_BID;
  (* RS_HS = "m_axi_in_47_B.ready" *)output m_axi_in_47_BREADY;
  (* RS_HS = "m_axi_in_47_B.data" *)input [1:0] m_axi_in_47_BRESP;
  (* RS_HS = "m_axi_in_47_B.valid" *)input m_axi_in_47_BVALID;
  (* RS_HS = "m_axi_in_47_R.data" *)input [255:0] m_axi_in_47_RDATA;
  (* RS_HS = "m_axi_in_47_R.data" *)input [0:0] m_axi_in_47_RID;
  (* RS_HS = "m_axi_in_47_R.data" *)input m_axi_in_47_RLAST;
  (* RS_HS = "m_axi_in_47_R.ready" *)output m_axi_in_47_RREADY;
  (* RS_HS = "m_axi_in_47_R.data" *)input [1:0] m_axi_in_47_RRESP;
  (* RS_HS = "m_axi_in_47_R.valid" *)input m_axi_in_47_RVALID;
  (* RS_HS = "m_axi_in_47_W.data" *)output [255:0] m_axi_in_47_WDATA;
  (* RS_HS = "m_axi_in_47_W.data" *)output m_axi_in_47_WLAST;
  (* RS_HS = "m_axi_in_47_W.ready" *)input m_axi_in_47_WREADY;
  (* RS_HS = "m_axi_in_47_W.data" *)output [31:0] m_axi_in_47_WSTRB;
  (* RS_HS = "m_axi_in_47_W.valid" *)output m_axi_in_47_WVALID;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [63:0] m_axi_in_48_ARADDR;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [1:0] m_axi_in_48_ARBURST;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [3:0] m_axi_in_48_ARCACHE;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [0:0] m_axi_in_48_ARID;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [7:0] m_axi_in_48_ARLEN;
  (* RS_HS = "m_axi_in_48_AR.data" *)output m_axi_in_48_ARLOCK;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [2:0] m_axi_in_48_ARPROT;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [3:0] m_axi_in_48_ARQOS;
  (* RS_HS = "m_axi_in_48_AR.ready" *)input m_axi_in_48_ARREADY;
  (* RS_HS = "m_axi_in_48_AR.data" *)output [2:0] m_axi_in_48_ARSIZE;
  (* RS_HS = "m_axi_in_48_AR.valid" *)output m_axi_in_48_ARVALID;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [63:0] m_axi_in_48_AWADDR;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [1:0] m_axi_in_48_AWBURST;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [3:0] m_axi_in_48_AWCACHE;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [0:0] m_axi_in_48_AWID;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [7:0] m_axi_in_48_AWLEN;
  (* RS_HS = "m_axi_in_48_AW.data" *)output m_axi_in_48_AWLOCK;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [2:0] m_axi_in_48_AWPROT;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [3:0] m_axi_in_48_AWQOS;
  (* RS_HS = "m_axi_in_48_AW.ready" *)input m_axi_in_48_AWREADY;
  (* RS_HS = "m_axi_in_48_AW.data" *)output [2:0] m_axi_in_48_AWSIZE;
  (* RS_HS = "m_axi_in_48_AW.valid" *)output m_axi_in_48_AWVALID;
  (* RS_HS = "m_axi_in_48_B.data" *)input [0:0] m_axi_in_48_BID;
  (* RS_HS = "m_axi_in_48_B.ready" *)output m_axi_in_48_BREADY;
  (* RS_HS = "m_axi_in_48_B.data" *)input [1:0] m_axi_in_48_BRESP;
  (* RS_HS = "m_axi_in_48_B.valid" *)input m_axi_in_48_BVALID;
  (* RS_HS = "m_axi_in_48_R.data" *)input [255:0] m_axi_in_48_RDATA;
  (* RS_HS = "m_axi_in_48_R.data" *)input [0:0] m_axi_in_48_RID;
  (* RS_HS = "m_axi_in_48_R.data" *)input m_axi_in_48_RLAST;
  (* RS_HS = "m_axi_in_48_R.ready" *)output m_axi_in_48_RREADY;
  (* RS_HS = "m_axi_in_48_R.data" *)input [1:0] m_axi_in_48_RRESP;
  (* RS_HS = "m_axi_in_48_R.valid" *)input m_axi_in_48_RVALID;
  (* RS_HS = "m_axi_in_48_W.data" *)output [255:0] m_axi_in_48_WDATA;
  (* RS_HS = "m_axi_in_48_W.data" *)output m_axi_in_48_WLAST;
  (* RS_HS = "m_axi_in_48_W.ready" *)input m_axi_in_48_WREADY;
  (* RS_HS = "m_axi_in_48_W.data" *)output [31:0] m_axi_in_48_WSTRB;
  (* RS_HS = "m_axi_in_48_W.valid" *)output m_axi_in_48_WVALID;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [63:0] m_axi_in_49_ARADDR;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [1:0] m_axi_in_49_ARBURST;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [3:0] m_axi_in_49_ARCACHE;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [0:0] m_axi_in_49_ARID;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [7:0] m_axi_in_49_ARLEN;
  (* RS_HS = "m_axi_in_49_AR.data" *)output m_axi_in_49_ARLOCK;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [2:0] m_axi_in_49_ARPROT;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [3:0] m_axi_in_49_ARQOS;
  (* RS_HS = "m_axi_in_49_AR.ready" *)input m_axi_in_49_ARREADY;
  (* RS_HS = "m_axi_in_49_AR.data" *)output [2:0] m_axi_in_49_ARSIZE;
  (* RS_HS = "m_axi_in_49_AR.valid" *)output m_axi_in_49_ARVALID;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [63:0] m_axi_in_49_AWADDR;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [1:0] m_axi_in_49_AWBURST;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [3:0] m_axi_in_49_AWCACHE;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [0:0] m_axi_in_49_AWID;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [7:0] m_axi_in_49_AWLEN;
  (* RS_HS = "m_axi_in_49_AW.data" *)output m_axi_in_49_AWLOCK;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [2:0] m_axi_in_49_AWPROT;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [3:0] m_axi_in_49_AWQOS;
  (* RS_HS = "m_axi_in_49_AW.ready" *)input m_axi_in_49_AWREADY;
  (* RS_HS = "m_axi_in_49_AW.data" *)output [2:0] m_axi_in_49_AWSIZE;
  (* RS_HS = "m_axi_in_49_AW.valid" *)output m_axi_in_49_AWVALID;
  (* RS_HS = "m_axi_in_49_B.data" *)input [0:0] m_axi_in_49_BID;
  (* RS_HS = "m_axi_in_49_B.ready" *)output m_axi_in_49_BREADY;
  (* RS_HS = "m_axi_in_49_B.data" *)input [1:0] m_axi_in_49_BRESP;
  (* RS_HS = "m_axi_in_49_B.valid" *)input m_axi_in_49_BVALID;
  (* RS_HS = "m_axi_in_49_R.data" *)input [255:0] m_axi_in_49_RDATA;
  (* RS_HS = "m_axi_in_49_R.data" *)input [0:0] m_axi_in_49_RID;
  (* RS_HS = "m_axi_in_49_R.data" *)input m_axi_in_49_RLAST;
  (* RS_HS = "m_axi_in_49_R.ready" *)output m_axi_in_49_RREADY;
  (* RS_HS = "m_axi_in_49_R.data" *)input [1:0] m_axi_in_49_RRESP;
  (* RS_HS = "m_axi_in_49_R.valid" *)input m_axi_in_49_RVALID;
  (* RS_HS = "m_axi_in_49_W.data" *)output [255:0] m_axi_in_49_WDATA;
  (* RS_HS = "m_axi_in_49_W.data" *)output m_axi_in_49_WLAST;
  (* RS_HS = "m_axi_in_49_W.ready" *)input m_axi_in_49_WREADY;
  (* RS_HS = "m_axi_in_49_W.data" *)output [31:0] m_axi_in_49_WSTRB;
  (* RS_HS = "m_axi_in_49_W.valid" *)output m_axi_in_49_WVALID;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [63:0] m_axi_in_5_ARADDR;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [1:0] m_axi_in_5_ARBURST;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [3:0] m_axi_in_5_ARCACHE;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [0:0] m_axi_in_5_ARID;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [7:0] m_axi_in_5_ARLEN;
  (* RS_HS = "m_axi_in_5_AR.data" *)output m_axi_in_5_ARLOCK;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [2:0] m_axi_in_5_ARPROT;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [3:0] m_axi_in_5_ARQOS;
  (* RS_HS = "m_axi_in_5_AR.ready" *)input m_axi_in_5_ARREADY;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [2:0] m_axi_in_5_ARSIZE;
  (* RS_HS = "m_axi_in_5_AR.valid" *)output m_axi_in_5_ARVALID;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [63:0] m_axi_in_5_AWADDR;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [1:0] m_axi_in_5_AWBURST;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [3:0] m_axi_in_5_AWCACHE;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [0:0] m_axi_in_5_AWID;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [7:0] m_axi_in_5_AWLEN;
  (* RS_HS = "m_axi_in_5_AW.data" *)output m_axi_in_5_AWLOCK;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [2:0] m_axi_in_5_AWPROT;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [3:0] m_axi_in_5_AWQOS;
  (* RS_HS = "m_axi_in_5_AW.ready" *)input m_axi_in_5_AWREADY;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [2:0] m_axi_in_5_AWSIZE;
  (* RS_HS = "m_axi_in_5_AW.valid" *)output m_axi_in_5_AWVALID;
  (* RS_HS = "m_axi_in_5_B.data" *)input [0:0] m_axi_in_5_BID;
  (* RS_HS = "m_axi_in_5_B.ready" *)output m_axi_in_5_BREADY;
  (* RS_HS = "m_axi_in_5_B.data" *)input [1:0] m_axi_in_5_BRESP;
  (* RS_HS = "m_axi_in_5_B.valid" *)input m_axi_in_5_BVALID;
  (* RS_HS = "m_axi_in_5_R.data" *)input [255:0] m_axi_in_5_RDATA;
  (* RS_HS = "m_axi_in_5_R.data" *)input [0:0] m_axi_in_5_RID;
  (* RS_HS = "m_axi_in_5_R.data" *)input m_axi_in_5_RLAST;
  (* RS_HS = "m_axi_in_5_R.ready" *)output m_axi_in_5_RREADY;
  (* RS_HS = "m_axi_in_5_R.data" *)input [1:0] m_axi_in_5_RRESP;
  (* RS_HS = "m_axi_in_5_R.valid" *)input m_axi_in_5_RVALID;
  (* RS_HS = "m_axi_in_5_W.data" *)output [255:0] m_axi_in_5_WDATA;
  (* RS_HS = "m_axi_in_5_W.data" *)output m_axi_in_5_WLAST;
  (* RS_HS = "m_axi_in_5_W.ready" *)input m_axi_in_5_WREADY;
  (* RS_HS = "m_axi_in_5_W.data" *)output [31:0] m_axi_in_5_WSTRB;
  (* RS_HS = "m_axi_in_5_W.valid" *)output m_axi_in_5_WVALID;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [63:0] m_axi_in_50_ARADDR;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [1:0] m_axi_in_50_ARBURST;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [3:0] m_axi_in_50_ARCACHE;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [0:0] m_axi_in_50_ARID;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [7:0] m_axi_in_50_ARLEN;
  (* RS_HS = "m_axi_in_50_AR.data" *)output m_axi_in_50_ARLOCK;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [2:0] m_axi_in_50_ARPROT;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [3:0] m_axi_in_50_ARQOS;
  (* RS_HS = "m_axi_in_50_AR.ready" *)input m_axi_in_50_ARREADY;
  (* RS_HS = "m_axi_in_50_AR.data" *)output [2:0] m_axi_in_50_ARSIZE;
  (* RS_HS = "m_axi_in_50_AR.valid" *)output m_axi_in_50_ARVALID;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [63:0] m_axi_in_50_AWADDR;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [1:0] m_axi_in_50_AWBURST;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [3:0] m_axi_in_50_AWCACHE;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [0:0] m_axi_in_50_AWID;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [7:0] m_axi_in_50_AWLEN;
  (* RS_HS = "m_axi_in_50_AW.data" *)output m_axi_in_50_AWLOCK;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [2:0] m_axi_in_50_AWPROT;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [3:0] m_axi_in_50_AWQOS;
  (* RS_HS = "m_axi_in_50_AW.ready" *)input m_axi_in_50_AWREADY;
  (* RS_HS = "m_axi_in_50_AW.data" *)output [2:0] m_axi_in_50_AWSIZE;
  (* RS_HS = "m_axi_in_50_AW.valid" *)output m_axi_in_50_AWVALID;
  (* RS_HS = "m_axi_in_50_B.data" *)input [0:0] m_axi_in_50_BID;
  (* RS_HS = "m_axi_in_50_B.ready" *)output m_axi_in_50_BREADY;
  (* RS_HS = "m_axi_in_50_B.data" *)input [1:0] m_axi_in_50_BRESP;
  (* RS_HS = "m_axi_in_50_B.valid" *)input m_axi_in_50_BVALID;
  (* RS_HS = "m_axi_in_50_R.data" *)input [255:0] m_axi_in_50_RDATA;
  (* RS_HS = "m_axi_in_50_R.data" *)input [0:0] m_axi_in_50_RID;
  (* RS_HS = "m_axi_in_50_R.data" *)input m_axi_in_50_RLAST;
  (* RS_HS = "m_axi_in_50_R.ready" *)output m_axi_in_50_RREADY;
  (* RS_HS = "m_axi_in_50_R.data" *)input [1:0] m_axi_in_50_RRESP;
  (* RS_HS = "m_axi_in_50_R.valid" *)input m_axi_in_50_RVALID;
  (* RS_HS = "m_axi_in_50_W.data" *)output [255:0] m_axi_in_50_WDATA;
  (* RS_HS = "m_axi_in_50_W.data" *)output m_axi_in_50_WLAST;
  (* RS_HS = "m_axi_in_50_W.ready" *)input m_axi_in_50_WREADY;
  (* RS_HS = "m_axi_in_50_W.data" *)output [31:0] m_axi_in_50_WSTRB;
  (* RS_HS = "m_axi_in_50_W.valid" *)output m_axi_in_50_WVALID;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [63:0] m_axi_in_51_ARADDR;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [1:0] m_axi_in_51_ARBURST;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [3:0] m_axi_in_51_ARCACHE;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [0:0] m_axi_in_51_ARID;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [7:0] m_axi_in_51_ARLEN;
  (* RS_HS = "m_axi_in_51_AR.data" *)output m_axi_in_51_ARLOCK;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [2:0] m_axi_in_51_ARPROT;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [3:0] m_axi_in_51_ARQOS;
  (* RS_HS = "m_axi_in_51_AR.ready" *)input m_axi_in_51_ARREADY;
  (* RS_HS = "m_axi_in_51_AR.data" *)output [2:0] m_axi_in_51_ARSIZE;
  (* RS_HS = "m_axi_in_51_AR.valid" *)output m_axi_in_51_ARVALID;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [63:0] m_axi_in_51_AWADDR;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [1:0] m_axi_in_51_AWBURST;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [3:0] m_axi_in_51_AWCACHE;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [0:0] m_axi_in_51_AWID;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [7:0] m_axi_in_51_AWLEN;
  (* RS_HS = "m_axi_in_51_AW.data" *)output m_axi_in_51_AWLOCK;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [2:0] m_axi_in_51_AWPROT;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [3:0] m_axi_in_51_AWQOS;
  (* RS_HS = "m_axi_in_51_AW.ready" *)input m_axi_in_51_AWREADY;
  (* RS_HS = "m_axi_in_51_AW.data" *)output [2:0] m_axi_in_51_AWSIZE;
  (* RS_HS = "m_axi_in_51_AW.valid" *)output m_axi_in_51_AWVALID;
  (* RS_HS = "m_axi_in_51_B.data" *)input [0:0] m_axi_in_51_BID;
  (* RS_HS = "m_axi_in_51_B.ready" *)output m_axi_in_51_BREADY;
  (* RS_HS = "m_axi_in_51_B.data" *)input [1:0] m_axi_in_51_BRESP;
  (* RS_HS = "m_axi_in_51_B.valid" *)input m_axi_in_51_BVALID;
  (* RS_HS = "m_axi_in_51_R.data" *)input [255:0] m_axi_in_51_RDATA;
  (* RS_HS = "m_axi_in_51_R.data" *)input [0:0] m_axi_in_51_RID;
  (* RS_HS = "m_axi_in_51_R.data" *)input m_axi_in_51_RLAST;
  (* RS_HS = "m_axi_in_51_R.ready" *)output m_axi_in_51_RREADY;
  (* RS_HS = "m_axi_in_51_R.data" *)input [1:0] m_axi_in_51_RRESP;
  (* RS_HS = "m_axi_in_51_R.valid" *)input m_axi_in_51_RVALID;
  (* RS_HS = "m_axi_in_51_W.data" *)output [255:0] m_axi_in_51_WDATA;
  (* RS_HS = "m_axi_in_51_W.data" *)output m_axi_in_51_WLAST;
  (* RS_HS = "m_axi_in_51_W.ready" *)input m_axi_in_51_WREADY;
  (* RS_HS = "m_axi_in_51_W.data" *)output [31:0] m_axi_in_51_WSTRB;
  (* RS_HS = "m_axi_in_51_W.valid" *)output m_axi_in_51_WVALID;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [63:0] m_axi_in_52_ARADDR;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [1:0] m_axi_in_52_ARBURST;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [3:0] m_axi_in_52_ARCACHE;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [0:0] m_axi_in_52_ARID;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [7:0] m_axi_in_52_ARLEN;
  (* RS_HS = "m_axi_in_52_AR.data" *)output m_axi_in_52_ARLOCK;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [2:0] m_axi_in_52_ARPROT;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [3:0] m_axi_in_52_ARQOS;
  (* RS_HS = "m_axi_in_52_AR.ready" *)input m_axi_in_52_ARREADY;
  (* RS_HS = "m_axi_in_52_AR.data" *)output [2:0] m_axi_in_52_ARSIZE;
  (* RS_HS = "m_axi_in_52_AR.valid" *)output m_axi_in_52_ARVALID;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [63:0] m_axi_in_52_AWADDR;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [1:0] m_axi_in_52_AWBURST;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [3:0] m_axi_in_52_AWCACHE;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [0:0] m_axi_in_52_AWID;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [7:0] m_axi_in_52_AWLEN;
  (* RS_HS = "m_axi_in_52_AW.data" *)output m_axi_in_52_AWLOCK;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [2:0] m_axi_in_52_AWPROT;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [3:0] m_axi_in_52_AWQOS;
  (* RS_HS = "m_axi_in_52_AW.ready" *)input m_axi_in_52_AWREADY;
  (* RS_HS = "m_axi_in_52_AW.data" *)output [2:0] m_axi_in_52_AWSIZE;
  (* RS_HS = "m_axi_in_52_AW.valid" *)output m_axi_in_52_AWVALID;
  (* RS_HS = "m_axi_in_52_B.data" *)input [0:0] m_axi_in_52_BID;
  (* RS_HS = "m_axi_in_52_B.ready" *)output m_axi_in_52_BREADY;
  (* RS_HS = "m_axi_in_52_B.data" *)input [1:0] m_axi_in_52_BRESP;
  (* RS_HS = "m_axi_in_52_B.valid" *)input m_axi_in_52_BVALID;
  (* RS_HS = "m_axi_in_52_R.data" *)input [255:0] m_axi_in_52_RDATA;
  (* RS_HS = "m_axi_in_52_R.data" *)input [0:0] m_axi_in_52_RID;
  (* RS_HS = "m_axi_in_52_R.data" *)input m_axi_in_52_RLAST;
  (* RS_HS = "m_axi_in_52_R.ready" *)output m_axi_in_52_RREADY;
  (* RS_HS = "m_axi_in_52_R.data" *)input [1:0] m_axi_in_52_RRESP;
  (* RS_HS = "m_axi_in_52_R.valid" *)input m_axi_in_52_RVALID;
  (* RS_HS = "m_axi_in_52_W.data" *)output [255:0] m_axi_in_52_WDATA;
  (* RS_HS = "m_axi_in_52_W.data" *)output m_axi_in_52_WLAST;
  (* RS_HS = "m_axi_in_52_W.ready" *)input m_axi_in_52_WREADY;
  (* RS_HS = "m_axi_in_52_W.data" *)output [31:0] m_axi_in_52_WSTRB;
  (* RS_HS = "m_axi_in_52_W.valid" *)output m_axi_in_52_WVALID;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [63:0] m_axi_in_53_ARADDR;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [1:0] m_axi_in_53_ARBURST;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [3:0] m_axi_in_53_ARCACHE;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [0:0] m_axi_in_53_ARID;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [7:0] m_axi_in_53_ARLEN;
  (* RS_HS = "m_axi_in_53_AR.data" *)output m_axi_in_53_ARLOCK;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [2:0] m_axi_in_53_ARPROT;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [3:0] m_axi_in_53_ARQOS;
  (* RS_HS = "m_axi_in_53_AR.ready" *)input m_axi_in_53_ARREADY;
  (* RS_HS = "m_axi_in_53_AR.data" *)output [2:0] m_axi_in_53_ARSIZE;
  (* RS_HS = "m_axi_in_53_AR.valid" *)output m_axi_in_53_ARVALID;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [63:0] m_axi_in_53_AWADDR;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [1:0] m_axi_in_53_AWBURST;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [3:0] m_axi_in_53_AWCACHE;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [0:0] m_axi_in_53_AWID;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [7:0] m_axi_in_53_AWLEN;
  (* RS_HS = "m_axi_in_53_AW.data" *)output m_axi_in_53_AWLOCK;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [2:0] m_axi_in_53_AWPROT;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [3:0] m_axi_in_53_AWQOS;
  (* RS_HS = "m_axi_in_53_AW.ready" *)input m_axi_in_53_AWREADY;
  (* RS_HS = "m_axi_in_53_AW.data" *)output [2:0] m_axi_in_53_AWSIZE;
  (* RS_HS = "m_axi_in_53_AW.valid" *)output m_axi_in_53_AWVALID;
  (* RS_HS = "m_axi_in_53_B.data" *)input [0:0] m_axi_in_53_BID;
  (* RS_HS = "m_axi_in_53_B.ready" *)output m_axi_in_53_BREADY;
  (* RS_HS = "m_axi_in_53_B.data" *)input [1:0] m_axi_in_53_BRESP;
  (* RS_HS = "m_axi_in_53_B.valid" *)input m_axi_in_53_BVALID;
  (* RS_HS = "m_axi_in_53_R.data" *)input [255:0] m_axi_in_53_RDATA;
  (* RS_HS = "m_axi_in_53_R.data" *)input [0:0] m_axi_in_53_RID;
  (* RS_HS = "m_axi_in_53_R.data" *)input m_axi_in_53_RLAST;
  (* RS_HS = "m_axi_in_53_R.ready" *)output m_axi_in_53_RREADY;
  (* RS_HS = "m_axi_in_53_R.data" *)input [1:0] m_axi_in_53_RRESP;
  (* RS_HS = "m_axi_in_53_R.valid" *)input m_axi_in_53_RVALID;
  (* RS_HS = "m_axi_in_53_W.data" *)output [255:0] m_axi_in_53_WDATA;
  (* RS_HS = "m_axi_in_53_W.data" *)output m_axi_in_53_WLAST;
  (* RS_HS = "m_axi_in_53_W.ready" *)input m_axi_in_53_WREADY;
  (* RS_HS = "m_axi_in_53_W.data" *)output [31:0] m_axi_in_53_WSTRB;
  (* RS_HS = "m_axi_in_53_W.valid" *)output m_axi_in_53_WVALID;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [63:0] m_axi_in_6_ARADDR;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [1:0] m_axi_in_6_ARBURST;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [3:0] m_axi_in_6_ARCACHE;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [0:0] m_axi_in_6_ARID;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [7:0] m_axi_in_6_ARLEN;
  (* RS_HS = "m_axi_in_6_AR.data" *)output m_axi_in_6_ARLOCK;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [2:0] m_axi_in_6_ARPROT;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [3:0] m_axi_in_6_ARQOS;
  (* RS_HS = "m_axi_in_6_AR.ready" *)input m_axi_in_6_ARREADY;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [2:0] m_axi_in_6_ARSIZE;
  (* RS_HS = "m_axi_in_6_AR.valid" *)output m_axi_in_6_ARVALID;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [63:0] m_axi_in_6_AWADDR;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [1:0] m_axi_in_6_AWBURST;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [3:0] m_axi_in_6_AWCACHE;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [0:0] m_axi_in_6_AWID;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [7:0] m_axi_in_6_AWLEN;
  (* RS_HS = "m_axi_in_6_AW.data" *)output m_axi_in_6_AWLOCK;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [2:0] m_axi_in_6_AWPROT;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [3:0] m_axi_in_6_AWQOS;
  (* RS_HS = "m_axi_in_6_AW.ready" *)input m_axi_in_6_AWREADY;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [2:0] m_axi_in_6_AWSIZE;
  (* RS_HS = "m_axi_in_6_AW.valid" *)output m_axi_in_6_AWVALID;
  (* RS_HS = "m_axi_in_6_B.data" *)input [0:0] m_axi_in_6_BID;
  (* RS_HS = "m_axi_in_6_B.ready" *)output m_axi_in_6_BREADY;
  (* RS_HS = "m_axi_in_6_B.data" *)input [1:0] m_axi_in_6_BRESP;
  (* RS_HS = "m_axi_in_6_B.valid" *)input m_axi_in_6_BVALID;
  (* RS_HS = "m_axi_in_6_R.data" *)input [255:0] m_axi_in_6_RDATA;
  (* RS_HS = "m_axi_in_6_R.data" *)input [0:0] m_axi_in_6_RID;
  (* RS_HS = "m_axi_in_6_R.data" *)input m_axi_in_6_RLAST;
  (* RS_HS = "m_axi_in_6_R.ready" *)output m_axi_in_6_RREADY;
  (* RS_HS = "m_axi_in_6_R.data" *)input [1:0] m_axi_in_6_RRESP;
  (* RS_HS = "m_axi_in_6_R.valid" *)input m_axi_in_6_RVALID;
  (* RS_HS = "m_axi_in_6_W.data" *)output [255:0] m_axi_in_6_WDATA;
  (* RS_HS = "m_axi_in_6_W.data" *)output m_axi_in_6_WLAST;
  (* RS_HS = "m_axi_in_6_W.ready" *)input m_axi_in_6_WREADY;
  (* RS_HS = "m_axi_in_6_W.data" *)output [31:0] m_axi_in_6_WSTRB;
  (* RS_HS = "m_axi_in_6_W.valid" *)output m_axi_in_6_WVALID;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [63:0] m_axi_in_7_ARADDR;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [1:0] m_axi_in_7_ARBURST;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [3:0] m_axi_in_7_ARCACHE;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [0:0] m_axi_in_7_ARID;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [7:0] m_axi_in_7_ARLEN;
  (* RS_HS = "m_axi_in_7_AR.data" *)output m_axi_in_7_ARLOCK;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [2:0] m_axi_in_7_ARPROT;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [3:0] m_axi_in_7_ARQOS;
  (* RS_HS = "m_axi_in_7_AR.ready" *)input m_axi_in_7_ARREADY;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [2:0] m_axi_in_7_ARSIZE;
  (* RS_HS = "m_axi_in_7_AR.valid" *)output m_axi_in_7_ARVALID;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [63:0] m_axi_in_7_AWADDR;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [1:0] m_axi_in_7_AWBURST;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [3:0] m_axi_in_7_AWCACHE;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [0:0] m_axi_in_7_AWID;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [7:0] m_axi_in_7_AWLEN;
  (* RS_HS = "m_axi_in_7_AW.data" *)output m_axi_in_7_AWLOCK;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [2:0] m_axi_in_7_AWPROT;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [3:0] m_axi_in_7_AWQOS;
  (* RS_HS = "m_axi_in_7_AW.ready" *)input m_axi_in_7_AWREADY;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [2:0] m_axi_in_7_AWSIZE;
  (* RS_HS = "m_axi_in_7_AW.valid" *)output m_axi_in_7_AWVALID;
  (* RS_HS = "m_axi_in_7_B.data" *)input [0:0] m_axi_in_7_BID;
  (* RS_HS = "m_axi_in_7_B.ready" *)output m_axi_in_7_BREADY;
  (* RS_HS = "m_axi_in_7_B.data" *)input [1:0] m_axi_in_7_BRESP;
  (* RS_HS = "m_axi_in_7_B.valid" *)input m_axi_in_7_BVALID;
  (* RS_HS = "m_axi_in_7_R.data" *)input [255:0] m_axi_in_7_RDATA;
  (* RS_HS = "m_axi_in_7_R.data" *)input [0:0] m_axi_in_7_RID;
  (* RS_HS = "m_axi_in_7_R.data" *)input m_axi_in_7_RLAST;
  (* RS_HS = "m_axi_in_7_R.ready" *)output m_axi_in_7_RREADY;
  (* RS_HS = "m_axi_in_7_R.data" *)input [1:0] m_axi_in_7_RRESP;
  (* RS_HS = "m_axi_in_7_R.valid" *)input m_axi_in_7_RVALID;
  (* RS_HS = "m_axi_in_7_W.data" *)output [255:0] m_axi_in_7_WDATA;
  (* RS_HS = "m_axi_in_7_W.data" *)output m_axi_in_7_WLAST;
  (* RS_HS = "m_axi_in_7_W.ready" *)input m_axi_in_7_WREADY;
  (* RS_HS = "m_axi_in_7_W.data" *)output [31:0] m_axi_in_7_WSTRB;
  (* RS_HS = "m_axi_in_7_W.valid" *)output m_axi_in_7_WVALID;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [63:0] m_axi_in_8_ARADDR;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [1:0] m_axi_in_8_ARBURST;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [3:0] m_axi_in_8_ARCACHE;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [0:0] m_axi_in_8_ARID;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [7:0] m_axi_in_8_ARLEN;
  (* RS_HS = "m_axi_in_8_AR.data" *)output m_axi_in_8_ARLOCK;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [2:0] m_axi_in_8_ARPROT;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [3:0] m_axi_in_8_ARQOS;
  (* RS_HS = "m_axi_in_8_AR.ready" *)input m_axi_in_8_ARREADY;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [2:0] m_axi_in_8_ARSIZE;
  (* RS_HS = "m_axi_in_8_AR.valid" *)output m_axi_in_8_ARVALID;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [63:0] m_axi_in_8_AWADDR;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [1:0] m_axi_in_8_AWBURST;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [3:0] m_axi_in_8_AWCACHE;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [0:0] m_axi_in_8_AWID;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [7:0] m_axi_in_8_AWLEN;
  (* RS_HS = "m_axi_in_8_AW.data" *)output m_axi_in_8_AWLOCK;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [2:0] m_axi_in_8_AWPROT;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [3:0] m_axi_in_8_AWQOS;
  (* RS_HS = "m_axi_in_8_AW.ready" *)input m_axi_in_8_AWREADY;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [2:0] m_axi_in_8_AWSIZE;
  (* RS_HS = "m_axi_in_8_AW.valid" *)output m_axi_in_8_AWVALID;
  (* RS_HS = "m_axi_in_8_B.data" *)input [0:0] m_axi_in_8_BID;
  (* RS_HS = "m_axi_in_8_B.ready" *)output m_axi_in_8_BREADY;
  (* RS_HS = "m_axi_in_8_B.data" *)input [1:0] m_axi_in_8_BRESP;
  (* RS_HS = "m_axi_in_8_B.valid" *)input m_axi_in_8_BVALID;
  (* RS_HS = "m_axi_in_8_R.data" *)input [255:0] m_axi_in_8_RDATA;
  (* RS_HS = "m_axi_in_8_R.data" *)input [0:0] m_axi_in_8_RID;
  (* RS_HS = "m_axi_in_8_R.data" *)input m_axi_in_8_RLAST;
  (* RS_HS = "m_axi_in_8_R.ready" *)output m_axi_in_8_RREADY;
  (* RS_HS = "m_axi_in_8_R.data" *)input [1:0] m_axi_in_8_RRESP;
  (* RS_HS = "m_axi_in_8_R.valid" *)input m_axi_in_8_RVALID;
  (* RS_HS = "m_axi_in_8_W.data" *)output [255:0] m_axi_in_8_WDATA;
  (* RS_HS = "m_axi_in_8_W.data" *)output m_axi_in_8_WLAST;
  (* RS_HS = "m_axi_in_8_W.ready" *)input m_axi_in_8_WREADY;
  (* RS_HS = "m_axi_in_8_W.data" *)output [31:0] m_axi_in_8_WSTRB;
  (* RS_HS = "m_axi_in_8_W.valid" *)output m_axi_in_8_WVALID;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [63:0] m_axi_in_9_ARADDR;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [1:0] m_axi_in_9_ARBURST;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [3:0] m_axi_in_9_ARCACHE;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [0:0] m_axi_in_9_ARID;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [7:0] m_axi_in_9_ARLEN;
  (* RS_HS = "m_axi_in_9_AR.data" *)output m_axi_in_9_ARLOCK;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [2:0] m_axi_in_9_ARPROT;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [3:0] m_axi_in_9_ARQOS;
  (* RS_HS = "m_axi_in_9_AR.ready" *)input m_axi_in_9_ARREADY;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [2:0] m_axi_in_9_ARSIZE;
  (* RS_HS = "m_axi_in_9_AR.valid" *)output m_axi_in_9_ARVALID;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [63:0] m_axi_in_9_AWADDR;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [1:0] m_axi_in_9_AWBURST;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [3:0] m_axi_in_9_AWCACHE;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [0:0] m_axi_in_9_AWID;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [7:0] m_axi_in_9_AWLEN;
  (* RS_HS = "m_axi_in_9_AW.data" *)output m_axi_in_9_AWLOCK;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [2:0] m_axi_in_9_AWPROT;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [3:0] m_axi_in_9_AWQOS;
  (* RS_HS = "m_axi_in_9_AW.ready" *)input m_axi_in_9_AWREADY;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [2:0] m_axi_in_9_AWSIZE;
  (* RS_HS = "m_axi_in_9_AW.valid" *)output m_axi_in_9_AWVALID;
  (* RS_HS = "m_axi_in_9_B.data" *)input [0:0] m_axi_in_9_BID;
  (* RS_HS = "m_axi_in_9_B.ready" *)output m_axi_in_9_BREADY;
  (* RS_HS = "m_axi_in_9_B.data" *)input [1:0] m_axi_in_9_BRESP;
  (* RS_HS = "m_axi_in_9_B.valid" *)input m_axi_in_9_BVALID;
  (* RS_HS = "m_axi_in_9_R.data" *)input [255:0] m_axi_in_9_RDATA;
  (* RS_HS = "m_axi_in_9_R.data" *)input [0:0] m_axi_in_9_RID;
  (* RS_HS = "m_axi_in_9_R.data" *)input m_axi_in_9_RLAST;
  (* RS_HS = "m_axi_in_9_R.ready" *)output m_axi_in_9_RREADY;
  (* RS_HS = "m_axi_in_9_R.data" *)input [1:0] m_axi_in_9_RRESP;
  (* RS_HS = "m_axi_in_9_R.valid" *)input m_axi_in_9_RVALID;
  (* RS_HS = "m_axi_in_9_W.data" *)output [255:0] m_axi_in_9_WDATA;
  (* RS_HS = "m_axi_in_9_W.data" *)output m_axi_in_9_WLAST;
  (* RS_HS = "m_axi_in_9_W.ready" *)input m_axi_in_9_WREADY;
  (* RS_HS = "m_axi_in_9_W.data" *)output [31:0] m_axi_in_9_WSTRB;
  (* RS_HS = "m_axi_in_9_W.valid" *)output m_axi_in_9_WVALID;
  wire ap_start;
  wire [63:0] in_0;
  wire [63:0] in_1;
  wire [63:0] in_2;
  wire [63:0] in_3;
  wire [63:0] in_4;
  wire [63:0] in_5;
  wire [63:0] in_6;
  wire [63:0] in_7;
  wire [63:0] in_8;
  wire [63:0] in_9;
  wire [63:0] in_10;
  wire [63:0] in_11;
  wire [63:0] in_12;
  wire [63:0] in_13;
  wire [63:0] in_14;
  wire [63:0] in_15;
  wire [63:0] in_16;
  wire [63:0] in_17;
  wire [63:0] in_18;
  wire [63:0] in_19;
  wire [63:0] in_20;
  wire [63:0] in_21;
  wire [63:0] in_22;
  wire [63:0] in_23;
  wire [63:0] in_24;
  wire [63:0] in_25;
  wire [63:0] in_26;
  wire [63:0] in_27;
  wire [63:0] in_28;
  wire [63:0] in_29;
  wire [63:0] in_30;
  wire [63:0] in_31;
  wire [63:0] in_32;
  wire [63:0] in_33;
  wire [63:0] in_34;
  wire [63:0] in_35;
  wire [63:0] in_36;
  wire [63:0] in_37;
  wire [63:0] in_38;
  wire [63:0] in_39;
  wire [63:0] in_40;
  wire [63:0] in_41;
  wire [63:0] in_42;
  wire [63:0] in_43;
  wire [63:0] in_44;
  wire [63:0] in_45;
  wire [63:0] in_46;
  wire [63:0] in_47;
  wire [63:0] in_48;
  wire [63:0] in_49;
  wire [63:0] in_50;
  wire [63:0] in_51;
  wire [63:0] in_52;
  wire [63:0] in_53;
  wire [63:0] L4_out_dist;
  wire [63:0] L4_out_id;
  wire [65:0] L1_out_dist_0__dout;
  wire L1_out_dist_0__empty_n;
  wire L1_out_dist_0__read;
  wire [65:0] L1_out_dist_0__din;
  wire L1_out_dist_0__full_n;
  wire L1_out_dist_0__write;
  wire [65:0] L1_out_dist_10__dout;
  wire L1_out_dist_10__empty_n;
  wire L1_out_dist_10__read;
  wire [65:0] L1_out_dist_10__din;
  wire L1_out_dist_10__full_n;
  wire L1_out_dist_10__write;
  wire [65:0] L1_out_dist_11__dout;
  wire L1_out_dist_11__empty_n;
  wire L1_out_dist_11__read;
  wire [65:0] L1_out_dist_11__din;
  wire L1_out_dist_11__full_n;
  wire L1_out_dist_11__write;
  wire [65:0] L1_out_dist_12__dout;
  wire L1_out_dist_12__empty_n;
  wire L1_out_dist_12__read;
  wire [65:0] L1_out_dist_12__din;
  wire L1_out_dist_12__full_n;
  wire L1_out_dist_12__write;
  wire [65:0] L1_out_dist_13__dout;
  wire L1_out_dist_13__empty_n;
  wire L1_out_dist_13__read;
  wire [65:0] L1_out_dist_13__din;
  wire L1_out_dist_13__full_n;
  wire L1_out_dist_13__write;
  wire [65:0] L1_out_dist_14__dout;
  wire L1_out_dist_14__empty_n;
  wire L1_out_dist_14__read;
  wire [65:0] L1_out_dist_14__din;
  wire L1_out_dist_14__full_n;
  wire L1_out_dist_14__write;
  wire [65:0] L1_out_dist_15__dout;
  wire L1_out_dist_15__empty_n;
  wire L1_out_dist_15__read;
  wire [65:0] L1_out_dist_15__din;
  wire L1_out_dist_15__full_n;
  wire L1_out_dist_15__write;
  wire [65:0] L1_out_dist_16__dout;
  wire L1_out_dist_16__empty_n;
  wire L1_out_dist_16__read;
  wire [65:0] L1_out_dist_16__din;
  wire L1_out_dist_16__full_n;
  wire L1_out_dist_16__write;
  wire [65:0] L1_out_dist_17__dout;
  wire L1_out_dist_17__empty_n;
  wire L1_out_dist_17__read;
  wire [65:0] L1_out_dist_17__din;
  wire L1_out_dist_17__full_n;
  wire L1_out_dist_17__write;
  wire [65:0] L1_out_dist_1__dout;
  wire L1_out_dist_1__empty_n;
  wire L1_out_dist_1__read;
  wire [65:0] L1_out_dist_1__din;
  wire L1_out_dist_1__full_n;
  wire L1_out_dist_1__write;
  wire [65:0] L1_out_dist_2__dout;
  wire L1_out_dist_2__empty_n;
  wire L1_out_dist_2__read;
  wire [65:0] L1_out_dist_2__din;
  wire L1_out_dist_2__full_n;
  wire L1_out_dist_2__write;
  wire [65:0] L1_out_dist_3__dout;
  wire L1_out_dist_3__empty_n;
  wire L1_out_dist_3__read;
  wire [65:0] L1_out_dist_3__din;
  wire L1_out_dist_3__full_n;
  wire L1_out_dist_3__write;
  wire [65:0] L1_out_dist_4__dout;
  wire L1_out_dist_4__empty_n;
  wire L1_out_dist_4__read;
  wire [65:0] L1_out_dist_4__din;
  wire L1_out_dist_4__full_n;
  wire L1_out_dist_4__write;
  wire [65:0] L1_out_dist_5__dout;
  wire L1_out_dist_5__empty_n;
  wire L1_out_dist_5__read;
  wire [65:0] L1_out_dist_5__din;
  wire L1_out_dist_5__full_n;
  wire L1_out_dist_5__write;
  wire [65:0] L1_out_dist_6__dout;
  wire L1_out_dist_6__empty_n;
  wire L1_out_dist_6__read;
  wire [65:0] L1_out_dist_6__din;
  wire L1_out_dist_6__full_n;
  wire L1_out_dist_6__write;
  wire [65:0] L1_out_dist_7__dout;
  wire L1_out_dist_7__empty_n;
  wire L1_out_dist_7__read;
  wire [65:0] L1_out_dist_7__din;
  wire L1_out_dist_7__full_n;
  wire L1_out_dist_7__write;
  wire [65:0] L1_out_dist_8__dout;
  wire L1_out_dist_8__empty_n;
  wire L1_out_dist_8__read;
  wire [65:0] L1_out_dist_8__din;
  wire L1_out_dist_8__full_n;
  wire L1_out_dist_8__write;
  wire [65:0] L1_out_dist_9__dout;
  wire L1_out_dist_9__empty_n;
  wire L1_out_dist_9__read;
  wire [65:0] L1_out_dist_9__din;
  wire L1_out_dist_9__full_n;
  wire L1_out_dist_9__write;
  wire [65:0] L1_out_id_0__dout;
  wire L1_out_id_0__empty_n;
  wire L1_out_id_0__read;
  wire [65:0] L1_out_id_0__din;
  wire L1_out_id_0__full_n;
  wire L1_out_id_0__write;
  wire [65:0] L1_out_id_10__dout;
  wire L1_out_id_10__empty_n;
  wire L1_out_id_10__read;
  wire [65:0] L1_out_id_10__din;
  wire L1_out_id_10__full_n;
  wire L1_out_id_10__write;
  wire [65:0] L1_out_id_11__dout;
  wire L1_out_id_11__empty_n;
  wire L1_out_id_11__read;
  wire [65:0] L1_out_id_11__din;
  wire L1_out_id_11__full_n;
  wire L1_out_id_11__write;
  wire [65:0] L1_out_id_12__dout;
  wire L1_out_id_12__empty_n;
  wire L1_out_id_12__read;
  wire [65:0] L1_out_id_12__din;
  wire L1_out_id_12__full_n;
  wire L1_out_id_12__write;
  wire [65:0] L1_out_id_13__dout;
  wire L1_out_id_13__empty_n;
  wire L1_out_id_13__read;
  wire [65:0] L1_out_id_13__din;
  wire L1_out_id_13__full_n;
  wire L1_out_id_13__write;
  wire [65:0] L1_out_id_14__dout;
  wire L1_out_id_14__empty_n;
  wire L1_out_id_14__read;
  wire [65:0] L1_out_id_14__din;
  wire L1_out_id_14__full_n;
  wire L1_out_id_14__write;
  wire [65:0] L1_out_id_15__dout;
  wire L1_out_id_15__empty_n;
  wire L1_out_id_15__read;
  wire [65:0] L1_out_id_15__din;
  wire L1_out_id_15__full_n;
  wire L1_out_id_15__write;
  wire [65:0] L1_out_id_16__dout;
  wire L1_out_id_16__empty_n;
  wire L1_out_id_16__read;
  wire [65:0] L1_out_id_16__din;
  wire L1_out_id_16__full_n;
  wire L1_out_id_16__write;
  wire [65:0] L1_out_id_17__dout;
  wire L1_out_id_17__empty_n;
  wire L1_out_id_17__read;
  wire [65:0] L1_out_id_17__din;
  wire L1_out_id_17__full_n;
  wire L1_out_id_17__write;
  wire [65:0] L1_out_id_1__dout;
  wire L1_out_id_1__empty_n;
  wire L1_out_id_1__read;
  wire [65:0] L1_out_id_1__din;
  wire L1_out_id_1__full_n;
  wire L1_out_id_1__write;
  wire [65:0] L1_out_id_2__dout;
  wire L1_out_id_2__empty_n;
  wire L1_out_id_2__read;
  wire [65:0] L1_out_id_2__din;
  wire L1_out_id_2__full_n;
  wire L1_out_id_2__write;
  wire [65:0] L1_out_id_3__dout;
  wire L1_out_id_3__empty_n;
  wire L1_out_id_3__read;
  wire [65:0] L1_out_id_3__din;
  wire L1_out_id_3__full_n;
  wire L1_out_id_3__write;
  wire [65:0] L1_out_id_4__dout;
  wire L1_out_id_4__empty_n;
  wire L1_out_id_4__read;
  wire [65:0] L1_out_id_4__din;
  wire L1_out_id_4__full_n;
  wire L1_out_id_4__write;
  wire [65:0] L1_out_id_5__dout;
  wire L1_out_id_5__empty_n;
  wire L1_out_id_5__read;
  wire [65:0] L1_out_id_5__din;
  wire L1_out_id_5__full_n;
  wire L1_out_id_5__write;
  wire [65:0] L1_out_id_6__dout;
  wire L1_out_id_6__empty_n;
  wire L1_out_id_6__read;
  wire [65:0] L1_out_id_6__din;
  wire L1_out_id_6__full_n;
  wire L1_out_id_6__write;
  wire [65:0] L1_out_id_7__dout;
  wire L1_out_id_7__empty_n;
  wire L1_out_id_7__read;
  wire [65:0] L1_out_id_7__din;
  wire L1_out_id_7__full_n;
  wire L1_out_id_7__write;
  wire [65:0] L1_out_id_8__dout;
  wire L1_out_id_8__empty_n;
  wire L1_out_id_8__read;
  wire [65:0] L1_out_id_8__din;
  wire L1_out_id_8__full_n;
  wire L1_out_id_8__write;
  wire [65:0] L1_out_id_9__dout;
  wire L1_out_id_9__empty_n;
  wire L1_out_id_9__read;
  wire [65:0] L1_out_id_9__din;
  wire L1_out_id_9__full_n;
  wire L1_out_id_9__write;
  wire [65:0] L2_out_dist0__dout;
  wire L2_out_dist0__empty_n;
  wire L2_out_dist0__read;
  wire [65:0] L2_out_dist0__din;
  wire L2_out_dist0__full_n;
  wire L2_out_dist0__write;
  wire [65:0] L2_out_dist1__dout;
  wire L2_out_dist1__empty_n;
  wire L2_out_dist1__read;
  wire [65:0] L2_out_dist1__din;
  wire L2_out_dist1__full_n;
  wire L2_out_dist1__write;
  wire [65:0] L2_out_dist2__dout;
  wire L2_out_dist2__empty_n;
  wire L2_out_dist2__read;
  wire [65:0] L2_out_dist2__din;
  wire L2_out_dist2__full_n;
  wire L2_out_dist2__write;
  wire [65:0] L2_out_dist3__dout;
  wire L2_out_dist3__empty_n;
  wire L2_out_dist3__read;
  wire [65:0] L2_out_dist3__din;
  wire L2_out_dist3__full_n;
  wire L2_out_dist3__write;
  wire [65:0] L2_out_dist4__dout;
  wire L2_out_dist4__empty_n;
  wire L2_out_dist4__read;
  wire [65:0] L2_out_dist4__din;
  wire L2_out_dist4__full_n;
  wire L2_out_dist4__write;
  wire [65:0] L2_out_dist5__dout;
  wire L2_out_dist5__empty_n;
  wire L2_out_dist5__read;
  wire [65:0] L2_out_dist5__din;
  wire L2_out_dist5__full_n;
  wire L2_out_dist5__write;
  wire [65:0] L2_out_id0__dout;
  wire L2_out_id0__empty_n;
  wire L2_out_id0__read;
  wire [65:0] L2_out_id0__din;
  wire L2_out_id0__full_n;
  wire L2_out_id0__write;
  wire [65:0] L2_out_id1__dout;
  wire L2_out_id1__empty_n;
  wire L2_out_id1__read;
  wire [65:0] L2_out_id1__din;
  wire L2_out_id1__full_n;
  wire L2_out_id1__write;
  wire [65:0] L2_out_id2__dout;
  wire L2_out_id2__empty_n;
  wire L2_out_id2__read;
  wire [65:0] L2_out_id2__din;
  wire L2_out_id2__full_n;
  wire L2_out_id2__write;
  wire [65:0] L2_out_id3__dout;
  wire L2_out_id3__empty_n;
  wire L2_out_id3__read;
  wire [65:0] L2_out_id3__din;
  wire L2_out_id3__full_n;
  wire L2_out_id3__write;
  wire [65:0] L2_out_id4__dout;
  wire L2_out_id4__empty_n;
  wire L2_out_id4__read;
  wire [65:0] L2_out_id4__din;
  wire L2_out_id4__full_n;
  wire L2_out_id4__write;
  wire [65:0] L2_out_id5__dout;
  wire L2_out_id5__empty_n;
  wire L2_out_id5__read;
  wire [65:0] L2_out_id5__din;
  wire L2_out_id5__full_n;
  wire L2_out_id5__write;
  wire [65:0] L3_out_dist0__dout;
  wire L3_out_dist0__empty_n;
  wire L3_out_dist0__read;
  wire [65:0] L3_out_dist0__din;
  wire L3_out_dist0__full_n;
  wire L3_out_dist0__write;
  wire [65:0] L3_out_dist1__dout;
  wire L3_out_dist1__empty_n;
  wire L3_out_dist1__read;
  wire [65:0] L3_out_dist1__din;
  wire L3_out_dist1__full_n;
  wire L3_out_dist1__write;
  wire [65:0] L3_out_id0__dout;
  wire L3_out_id0__empty_n;
  wire L3_out_id0__read;
  wire [65:0] L3_out_id0__din;
  wire L3_out_id0__full_n;
  wire L3_out_id0__write;
  wire [65:0] L3_out_id1__dout;
  wire L3_out_id1__empty_n;
  wire L3_out_id1__read;
  wire [65:0] L3_out_id1__din;
  wire L3_out_id1__full_n;
  wire L3_out_id1__write;
  wire [65:0] out_dist_0__dout;
  wire out_dist_0__empty_n;
  wire out_dist_0__read;
  wire [65:0] out_dist_0__din;
  wire out_dist_0__full_n;
  wire out_dist_0__write;
  wire [65:0] out_dist_10__dout;
  wire out_dist_10__empty_n;
  wire out_dist_10__read;
  wire [65:0] out_dist_10__din;
  wire out_dist_10__full_n;
  wire out_dist_10__write;
  wire [65:0] out_dist_11__dout;
  wire out_dist_11__empty_n;
  wire out_dist_11__read;
  wire [65:0] out_dist_11__din;
  wire out_dist_11__full_n;
  wire out_dist_11__write;
  wire [65:0] out_dist_12__dout;
  wire out_dist_12__empty_n;
  wire out_dist_12__read;
  wire [65:0] out_dist_12__din;
  wire out_dist_12__full_n;
  wire out_dist_12__write;
  wire [65:0] out_dist_13__dout;
  wire out_dist_13__empty_n;
  wire out_dist_13__read;
  wire [65:0] out_dist_13__din;
  wire out_dist_13__full_n;
  wire out_dist_13__write;
  wire [65:0] out_dist_14__dout;
  wire out_dist_14__empty_n;
  wire out_dist_14__read;
  wire [65:0] out_dist_14__din;
  wire out_dist_14__full_n;
  wire out_dist_14__write;
  wire [65:0] out_dist_15__dout;
  wire out_dist_15__empty_n;
  wire out_dist_15__read;
  wire [65:0] out_dist_15__din;
  wire out_dist_15__full_n;
  wire out_dist_15__write;
  wire [65:0] out_dist_16__dout;
  wire out_dist_16__empty_n;
  wire out_dist_16__read;
  wire [65:0] out_dist_16__din;
  wire out_dist_16__full_n;
  wire out_dist_16__write;
  wire [65:0] out_dist_17__dout;
  wire out_dist_17__empty_n;
  wire out_dist_17__read;
  wire [65:0] out_dist_17__din;
  wire out_dist_17__full_n;
  wire out_dist_17__write;
  wire [65:0] out_dist_18__dout;
  wire out_dist_18__empty_n;
  wire out_dist_18__read;
  wire [65:0] out_dist_18__din;
  wire out_dist_18__full_n;
  wire out_dist_18__write;
  wire [65:0] out_dist_19__dout;
  wire out_dist_19__empty_n;
  wire out_dist_19__read;
  wire [65:0] out_dist_19__din;
  wire out_dist_19__full_n;
  wire out_dist_19__write;
  wire [65:0] out_dist_1__dout;
  wire out_dist_1__empty_n;
  wire out_dist_1__read;
  wire [65:0] out_dist_1__din;
  wire out_dist_1__full_n;
  wire out_dist_1__write;
  wire [65:0] out_dist_20__dout;
  wire out_dist_20__empty_n;
  wire out_dist_20__read;
  wire [65:0] out_dist_20__din;
  wire out_dist_20__full_n;
  wire out_dist_20__write;
  wire [65:0] out_dist_21__dout;
  wire out_dist_21__empty_n;
  wire out_dist_21__read;
  wire [65:0] out_dist_21__din;
  wire out_dist_21__full_n;
  wire out_dist_21__write;
  wire [65:0] out_dist_22__dout;
  wire out_dist_22__empty_n;
  wire out_dist_22__read;
  wire [65:0] out_dist_22__din;
  wire out_dist_22__full_n;
  wire out_dist_22__write;
  wire [65:0] out_dist_23__dout;
  wire out_dist_23__empty_n;
  wire out_dist_23__read;
  wire [65:0] out_dist_23__din;
  wire out_dist_23__full_n;
  wire out_dist_23__write;
  wire [65:0] out_dist_24__dout;
  wire out_dist_24__empty_n;
  wire out_dist_24__read;
  wire [65:0] out_dist_24__din;
  wire out_dist_24__full_n;
  wire out_dist_24__write;
  wire [65:0] out_dist_25__dout;
  wire out_dist_25__empty_n;
  wire out_dist_25__read;
  wire [65:0] out_dist_25__din;
  wire out_dist_25__full_n;
  wire out_dist_25__write;
  wire [65:0] out_dist_26__dout;
  wire out_dist_26__empty_n;
  wire out_dist_26__read;
  wire [65:0] out_dist_26__din;
  wire out_dist_26__full_n;
  wire out_dist_26__write;
  wire [65:0] out_dist_27__dout;
  wire out_dist_27__empty_n;
  wire out_dist_27__read;
  wire [65:0] out_dist_27__din;
  wire out_dist_27__full_n;
  wire out_dist_27__write;
  wire [65:0] out_dist_28__dout;
  wire out_dist_28__empty_n;
  wire out_dist_28__read;
  wire [65:0] out_dist_28__din;
  wire out_dist_28__full_n;
  wire out_dist_28__write;
  wire [65:0] out_dist_29__dout;
  wire out_dist_29__empty_n;
  wire out_dist_29__read;
  wire [65:0] out_dist_29__din;
  wire out_dist_29__full_n;
  wire out_dist_29__write;
  wire [65:0] out_dist_2__dout;
  wire out_dist_2__empty_n;
  wire out_dist_2__read;
  wire [65:0] out_dist_2__din;
  wire out_dist_2__full_n;
  wire out_dist_2__write;
  wire [65:0] out_dist_30__dout;
  wire out_dist_30__empty_n;
  wire out_dist_30__read;
  wire [65:0] out_dist_30__din;
  wire out_dist_30__full_n;
  wire out_dist_30__write;
  wire [65:0] out_dist_31__dout;
  wire out_dist_31__empty_n;
  wire out_dist_31__read;
  wire [65:0] out_dist_31__din;
  wire out_dist_31__full_n;
  wire out_dist_31__write;
  wire [65:0] out_dist_32__dout;
  wire out_dist_32__empty_n;
  wire out_dist_32__read;
  wire [65:0] out_dist_32__din;
  wire out_dist_32__full_n;
  wire out_dist_32__write;
  wire [65:0] out_dist_33__dout;
  wire out_dist_33__empty_n;
  wire out_dist_33__read;
  wire [65:0] out_dist_33__din;
  wire out_dist_33__full_n;
  wire out_dist_33__write;
  wire [65:0] out_dist_34__dout;
  wire out_dist_34__empty_n;
  wire out_dist_34__read;
  wire [65:0] out_dist_34__din;
  wire out_dist_34__full_n;
  wire out_dist_34__write;
  wire [65:0] out_dist_35__dout;
  wire out_dist_35__empty_n;
  wire out_dist_35__read;
  wire [65:0] out_dist_35__din;
  wire out_dist_35__full_n;
  wire out_dist_35__write;
  wire [65:0] out_dist_36__dout;
  wire out_dist_36__empty_n;
  wire out_dist_36__read;
  wire [65:0] out_dist_36__din;
  wire out_dist_36__full_n;
  wire out_dist_36__write;
  wire [65:0] out_dist_37__dout;
  wire out_dist_37__empty_n;
  wire out_dist_37__read;
  wire [65:0] out_dist_37__din;
  wire out_dist_37__full_n;
  wire out_dist_37__write;
  wire [65:0] out_dist_38__dout;
  wire out_dist_38__empty_n;
  wire out_dist_38__read;
  wire [65:0] out_dist_38__din;
  wire out_dist_38__full_n;
  wire out_dist_38__write;
  wire [65:0] out_dist_39__dout;
  wire out_dist_39__empty_n;
  wire out_dist_39__read;
  wire [65:0] out_dist_39__din;
  wire out_dist_39__full_n;
  wire out_dist_39__write;
  wire [65:0] out_dist_3__dout;
  wire out_dist_3__empty_n;
  wire out_dist_3__read;
  wire [65:0] out_dist_3__din;
  wire out_dist_3__full_n;
  wire out_dist_3__write;
  wire [65:0] out_dist_40__dout;
  wire out_dist_40__empty_n;
  wire out_dist_40__read;
  wire [65:0] out_dist_40__din;
  wire out_dist_40__full_n;
  wire out_dist_40__write;
  wire [65:0] out_dist_41__dout;
  wire out_dist_41__empty_n;
  wire out_dist_41__read;
  wire [65:0] out_dist_41__din;
  wire out_dist_41__full_n;
  wire out_dist_41__write;
  wire [65:0] out_dist_42__dout;
  wire out_dist_42__empty_n;
  wire out_dist_42__read;
  wire [65:0] out_dist_42__din;
  wire out_dist_42__full_n;
  wire out_dist_42__write;
  wire [65:0] out_dist_43__dout;
  wire out_dist_43__empty_n;
  wire out_dist_43__read;
  wire [65:0] out_dist_43__din;
  wire out_dist_43__full_n;
  wire out_dist_43__write;
  wire [65:0] out_dist_44__dout;
  wire out_dist_44__empty_n;
  wire out_dist_44__read;
  wire [65:0] out_dist_44__din;
  wire out_dist_44__full_n;
  wire out_dist_44__write;
  wire [65:0] out_dist_45__dout;
  wire out_dist_45__empty_n;
  wire out_dist_45__read;
  wire [65:0] out_dist_45__din;
  wire out_dist_45__full_n;
  wire out_dist_45__write;
  wire [65:0] out_dist_46__dout;
  wire out_dist_46__empty_n;
  wire out_dist_46__read;
  wire [65:0] out_dist_46__din;
  wire out_dist_46__full_n;
  wire out_dist_46__write;
  wire [65:0] out_dist_47__dout;
  wire out_dist_47__empty_n;
  wire out_dist_47__read;
  wire [65:0] out_dist_47__din;
  wire out_dist_47__full_n;
  wire out_dist_47__write;
  wire [65:0] out_dist_48__dout;
  wire out_dist_48__empty_n;
  wire out_dist_48__read;
  wire [65:0] out_dist_48__din;
  wire out_dist_48__full_n;
  wire out_dist_48__write;
  wire [65:0] out_dist_49__dout;
  wire out_dist_49__empty_n;
  wire out_dist_49__read;
  wire [65:0] out_dist_49__din;
  wire out_dist_49__full_n;
  wire out_dist_49__write;
  wire [65:0] out_dist_4__dout;
  wire out_dist_4__empty_n;
  wire out_dist_4__read;
  wire [65:0] out_dist_4__din;
  wire out_dist_4__full_n;
  wire out_dist_4__write;
  wire [65:0] out_dist_50__dout;
  wire out_dist_50__empty_n;
  wire out_dist_50__read;
  wire [65:0] out_dist_50__din;
  wire out_dist_50__full_n;
  wire out_dist_50__write;
  wire [65:0] out_dist_51__dout;
  wire out_dist_51__empty_n;
  wire out_dist_51__read;
  wire [65:0] out_dist_51__din;
  wire out_dist_51__full_n;
  wire out_dist_51__write;
  wire [65:0] out_dist_52__dout;
  wire out_dist_52__empty_n;
  wire out_dist_52__read;
  wire [65:0] out_dist_52__din;
  wire out_dist_52__full_n;
  wire out_dist_52__write;
  wire [65:0] out_dist_53__dout;
  wire out_dist_53__empty_n;
  wire out_dist_53__read;
  wire [65:0] out_dist_53__din;
  wire out_dist_53__full_n;
  wire out_dist_53__write;
  wire [65:0] out_dist_5__dout;
  wire out_dist_5__empty_n;
  wire out_dist_5__read;
  wire [65:0] out_dist_5__din;
  wire out_dist_5__full_n;
  wire out_dist_5__write;
  wire [65:0] out_dist_6__dout;
  wire out_dist_6__empty_n;
  wire out_dist_6__read;
  wire [65:0] out_dist_6__din;
  wire out_dist_6__full_n;
  wire out_dist_6__write;
  wire [65:0] out_dist_7__dout;
  wire out_dist_7__empty_n;
  wire out_dist_7__read;
  wire [65:0] out_dist_7__din;
  wire out_dist_7__full_n;
  wire out_dist_7__write;
  wire [65:0] out_dist_8__dout;
  wire out_dist_8__empty_n;
  wire out_dist_8__read;
  wire [65:0] out_dist_8__din;
  wire out_dist_8__full_n;
  wire out_dist_8__write;
  wire [65:0] out_dist_9__dout;
  wire out_dist_9__empty_n;
  wire out_dist_9__read;
  wire [65:0] out_dist_9__din;
  wire out_dist_9__full_n;
  wire out_dist_9__write;
  wire [65:0] out_id_0__dout;
  wire out_id_0__empty_n;
  wire out_id_0__read;
  wire [65:0] out_id_0__din;
  wire out_id_0__full_n;
  wire out_id_0__write;
  wire [65:0] out_id_10__dout;
  wire out_id_10__empty_n;
  wire out_id_10__read;
  wire [65:0] out_id_10__din;
  wire out_id_10__full_n;
  wire out_id_10__write;
  wire [65:0] out_id_11__dout;
  wire out_id_11__empty_n;
  wire out_id_11__read;
  wire [65:0] out_id_11__din;
  wire out_id_11__full_n;
  wire out_id_11__write;
  wire [65:0] out_id_12__dout;
  wire out_id_12__empty_n;
  wire out_id_12__read;
  wire [65:0] out_id_12__din;
  wire out_id_12__full_n;
  wire out_id_12__write;
  wire [65:0] out_id_13__dout;
  wire out_id_13__empty_n;
  wire out_id_13__read;
  wire [65:0] out_id_13__din;
  wire out_id_13__full_n;
  wire out_id_13__write;
  wire [65:0] out_id_14__dout;
  wire out_id_14__empty_n;
  wire out_id_14__read;
  wire [65:0] out_id_14__din;
  wire out_id_14__full_n;
  wire out_id_14__write;
  wire [65:0] out_id_15__dout;
  wire out_id_15__empty_n;
  wire out_id_15__read;
  wire [65:0] out_id_15__din;
  wire out_id_15__full_n;
  wire out_id_15__write;
  wire [65:0] out_id_16__dout;
  wire out_id_16__empty_n;
  wire out_id_16__read;
  wire [65:0] out_id_16__din;
  wire out_id_16__full_n;
  wire out_id_16__write;
  wire [65:0] out_id_17__dout;
  wire out_id_17__empty_n;
  wire out_id_17__read;
  wire [65:0] out_id_17__din;
  wire out_id_17__full_n;
  wire out_id_17__write;
  wire [65:0] out_id_18__dout;
  wire out_id_18__empty_n;
  wire out_id_18__read;
  wire [65:0] out_id_18__din;
  wire out_id_18__full_n;
  wire out_id_18__write;
  wire [65:0] out_id_19__dout;
  wire out_id_19__empty_n;
  wire out_id_19__read;
  wire [65:0] out_id_19__din;
  wire out_id_19__full_n;
  wire out_id_19__write;
  wire [65:0] out_id_1__dout;
  wire out_id_1__empty_n;
  wire out_id_1__read;
  wire [65:0] out_id_1__din;
  wire out_id_1__full_n;
  wire out_id_1__write;
  wire [65:0] out_id_20__dout;
  wire out_id_20__empty_n;
  wire out_id_20__read;
  wire [65:0] out_id_20__din;
  wire out_id_20__full_n;
  wire out_id_20__write;
  wire [65:0] out_id_21__dout;
  wire out_id_21__empty_n;
  wire out_id_21__read;
  wire [65:0] out_id_21__din;
  wire out_id_21__full_n;
  wire out_id_21__write;
  wire [65:0] out_id_22__dout;
  wire out_id_22__empty_n;
  wire out_id_22__read;
  wire [65:0] out_id_22__din;
  wire out_id_22__full_n;
  wire out_id_22__write;
  wire [65:0] out_id_23__dout;
  wire out_id_23__empty_n;
  wire out_id_23__read;
  wire [65:0] out_id_23__din;
  wire out_id_23__full_n;
  wire out_id_23__write;
  wire [65:0] out_id_24__dout;
  wire out_id_24__empty_n;
  wire out_id_24__read;
  wire [65:0] out_id_24__din;
  wire out_id_24__full_n;
  wire out_id_24__write;
  wire [65:0] out_id_25__dout;
  wire out_id_25__empty_n;
  wire out_id_25__read;
  wire [65:0] out_id_25__din;
  wire out_id_25__full_n;
  wire out_id_25__write;
  wire [65:0] out_id_26__dout;
  wire out_id_26__empty_n;
  wire out_id_26__read;
  wire [65:0] out_id_26__din;
  wire out_id_26__full_n;
  wire out_id_26__write;
  wire [65:0] out_id_27__dout;
  wire out_id_27__empty_n;
  wire out_id_27__read;
  wire [65:0] out_id_27__din;
  wire out_id_27__full_n;
  wire out_id_27__write;
  wire [65:0] out_id_28__dout;
  wire out_id_28__empty_n;
  wire out_id_28__read;
  wire [65:0] out_id_28__din;
  wire out_id_28__full_n;
  wire out_id_28__write;
  wire [65:0] out_id_29__dout;
  wire out_id_29__empty_n;
  wire out_id_29__read;
  wire [65:0] out_id_29__din;
  wire out_id_29__full_n;
  wire out_id_29__write;
  wire [65:0] out_id_2__dout;
  wire out_id_2__empty_n;
  wire out_id_2__read;
  wire [65:0] out_id_2__din;
  wire out_id_2__full_n;
  wire out_id_2__write;
  wire [65:0] out_id_30__dout;
  wire out_id_30__empty_n;
  wire out_id_30__read;
  wire [65:0] out_id_30__din;
  wire out_id_30__full_n;
  wire out_id_30__write;
  wire [65:0] out_id_31__dout;
  wire out_id_31__empty_n;
  wire out_id_31__read;
  wire [65:0] out_id_31__din;
  wire out_id_31__full_n;
  wire out_id_31__write;
  wire [65:0] out_id_32__dout;
  wire out_id_32__empty_n;
  wire out_id_32__read;
  wire [65:0] out_id_32__din;
  wire out_id_32__full_n;
  wire out_id_32__write;
  wire [65:0] out_id_33__dout;
  wire out_id_33__empty_n;
  wire out_id_33__read;
  wire [65:0] out_id_33__din;
  wire out_id_33__full_n;
  wire out_id_33__write;
  wire [65:0] out_id_34__dout;
  wire out_id_34__empty_n;
  wire out_id_34__read;
  wire [65:0] out_id_34__din;
  wire out_id_34__full_n;
  wire out_id_34__write;
  wire [65:0] out_id_35__dout;
  wire out_id_35__empty_n;
  wire out_id_35__read;
  wire [65:0] out_id_35__din;
  wire out_id_35__full_n;
  wire out_id_35__write;
  wire [65:0] out_id_36__dout;
  wire out_id_36__empty_n;
  wire out_id_36__read;
  wire [65:0] out_id_36__din;
  wire out_id_36__full_n;
  wire out_id_36__write;
  wire [65:0] out_id_37__dout;
  wire out_id_37__empty_n;
  wire out_id_37__read;
  wire [65:0] out_id_37__din;
  wire out_id_37__full_n;
  wire out_id_37__write;
  wire [65:0] out_id_38__dout;
  wire out_id_38__empty_n;
  wire out_id_38__read;
  wire [65:0] out_id_38__din;
  wire out_id_38__full_n;
  wire out_id_38__write;
  wire [65:0] out_id_39__dout;
  wire out_id_39__empty_n;
  wire out_id_39__read;
  wire [65:0] out_id_39__din;
  wire out_id_39__full_n;
  wire out_id_39__write;
  wire [65:0] out_id_3__dout;
  wire out_id_3__empty_n;
  wire out_id_3__read;
  wire [65:0] out_id_3__din;
  wire out_id_3__full_n;
  wire out_id_3__write;
  wire [65:0] out_id_40__dout;
  wire out_id_40__empty_n;
  wire out_id_40__read;
  wire [65:0] out_id_40__din;
  wire out_id_40__full_n;
  wire out_id_40__write;
  wire [65:0] out_id_41__dout;
  wire out_id_41__empty_n;
  wire out_id_41__read;
  wire [65:0] out_id_41__din;
  wire out_id_41__full_n;
  wire out_id_41__write;
  wire [65:0] out_id_42__dout;
  wire out_id_42__empty_n;
  wire out_id_42__read;
  wire [65:0] out_id_42__din;
  wire out_id_42__full_n;
  wire out_id_42__write;
  wire [65:0] out_id_43__dout;
  wire out_id_43__empty_n;
  wire out_id_43__read;
  wire [65:0] out_id_43__din;
  wire out_id_43__full_n;
  wire out_id_43__write;
  wire [65:0] out_id_44__dout;
  wire out_id_44__empty_n;
  wire out_id_44__read;
  wire [65:0] out_id_44__din;
  wire out_id_44__full_n;
  wire out_id_44__write;
  wire [65:0] out_id_45__dout;
  wire out_id_45__empty_n;
  wire out_id_45__read;
  wire [65:0] out_id_45__din;
  wire out_id_45__full_n;
  wire out_id_45__write;
  wire [65:0] out_id_46__dout;
  wire out_id_46__empty_n;
  wire out_id_46__read;
  wire [65:0] out_id_46__din;
  wire out_id_46__full_n;
  wire out_id_46__write;
  wire [65:0] out_id_47__dout;
  wire out_id_47__empty_n;
  wire out_id_47__read;
  wire [65:0] out_id_47__din;
  wire out_id_47__full_n;
  wire out_id_47__write;
  wire [65:0] out_id_48__dout;
  wire out_id_48__empty_n;
  wire out_id_48__read;
  wire [65:0] out_id_48__din;
  wire out_id_48__full_n;
  wire out_id_48__write;
  wire [65:0] out_id_49__dout;
  wire out_id_49__empty_n;
  wire out_id_49__read;
  wire [65:0] out_id_49__din;
  wire out_id_49__full_n;
  wire out_id_49__write;
  wire [65:0] out_id_4__dout;
  wire out_id_4__empty_n;
  wire out_id_4__read;
  wire [65:0] out_id_4__din;
  wire out_id_4__full_n;
  wire out_id_4__write;
  wire [65:0] out_id_50__dout;
  wire out_id_50__empty_n;
  wire out_id_50__read;
  wire [65:0] out_id_50__din;
  wire out_id_50__full_n;
  wire out_id_50__write;
  wire [65:0] out_id_51__dout;
  wire out_id_51__empty_n;
  wire out_id_51__read;
  wire [65:0] out_id_51__din;
  wire out_id_51__full_n;
  wire out_id_51__write;
  wire [65:0] out_id_52__dout;
  wire out_id_52__empty_n;
  wire out_id_52__read;
  wire [65:0] out_id_52__din;
  wire out_id_52__full_n;
  wire out_id_52__write;
  wire [65:0] out_id_53__dout;
  wire out_id_53__empty_n;
  wire out_id_53__read;
  wire [65:0] out_id_53__din;
  wire out_id_53__full_n;
  wire out_id_53__write;
  wire [65:0] out_id_5__dout;
  wire out_id_5__empty_n;
  wire out_id_5__read;
  wire [65:0] out_id_5__din;
  wire out_id_5__full_n;
  wire out_id_5__write;
  wire [65:0] out_id_6__dout;
  wire out_id_6__empty_n;
  wire out_id_6__read;
  wire [65:0] out_id_6__din;
  wire out_id_6__full_n;
  wire out_id_6__write;
  wire [65:0] out_id_7__dout;
  wire out_id_7__empty_n;
  wire out_id_7__read;
  wire [65:0] out_id_7__din;
  wire out_id_7__full_n;
  wire out_id_7__write;
  wire [65:0] out_id_8__dout;
  wire out_id_8__empty_n;
  wire out_id_8__read;
  wire [65:0] out_id_8__din;
  wire out_id_8__full_n;
  wire out_id_8__write;
  wire [65:0] out_id_9__dout;
  wire out_id_9__empty_n;
  wire out_id_9__read;
  wire [65:0] out_id_9__din;
  wire out_id_9__full_n;
  wire out_id_9__write;
  wire krnl_globalSort_L1_L2_0__ap_start;
  wire krnl_globalSort_L1_L2_0__ap_ready;
  wire krnl_globalSort_L1_L2_0__ap_done;
  wire krnl_globalSort_L1_L2_0__ap_idle;
  wire krnl_globalSort_L1_L2_1__ap_start;
  wire krnl_globalSort_L1_L2_1__ap_ready;
  wire krnl_globalSort_L1_L2_1__ap_done;
  wire krnl_globalSort_L1_L2_1__ap_idle;
  wire krnl_globalSort_L1_L2_2__ap_start;
  wire krnl_globalSort_L1_L2_2__ap_ready;
  wire krnl_globalSort_L1_L2_2__ap_done;
  wire krnl_globalSort_L1_L2_2__ap_idle;
  wire krnl_globalSort_L1_L2_3__ap_start;
  wire krnl_globalSort_L1_L2_3__ap_ready;
  wire krnl_globalSort_L1_L2_3__ap_done;
  wire krnl_globalSort_L1_L2_3__ap_idle;
  wire krnl_globalSort_L1_L2_4__ap_start;
  wire krnl_globalSort_L1_L2_4__ap_ready;
  wire krnl_globalSort_L1_L2_4__ap_done;
  wire krnl_globalSort_L1_L2_4__ap_idle;
  wire krnl_globalSort_L1_L2_5__ap_start;
  wire krnl_globalSort_L1_L2_5__ap_ready;
  wire krnl_globalSort_L1_L2_5__ap_done;
  wire krnl_globalSort_L1_L2_5__ap_idle;
  wire krnl_globalSort_L1_L2_6__ap_start;
  wire krnl_globalSort_L1_L2_6__ap_ready;
  wire krnl_globalSort_L1_L2_6__ap_done;
  wire krnl_globalSort_L1_L2_6__ap_idle;
  wire krnl_globalSort_L1_L2_7__ap_start;
  wire krnl_globalSort_L1_L2_7__ap_ready;
  wire krnl_globalSort_L1_L2_7__ap_done;
  wire krnl_globalSort_L1_L2_7__ap_idle;
  wire krnl_globalSort_L1_L2_8__ap_start;
  wire krnl_globalSort_L1_L2_8__ap_ready;
  wire krnl_globalSort_L1_L2_8__ap_done;
  wire krnl_globalSort_L1_L2_8__ap_idle;
  wire krnl_globalSort_L1_L2_9__ap_start;
  wire krnl_globalSort_L1_L2_9__ap_ready;
  wire krnl_globalSort_L1_L2_9__ap_done;
  wire krnl_globalSort_L1_L2_9__ap_idle;
  wire krnl_globalSort_L1_L2_10__ap_start;
  wire krnl_globalSort_L1_L2_10__ap_ready;
  wire krnl_globalSort_L1_L2_10__ap_done;
  wire krnl_globalSort_L1_L2_10__ap_idle;
  wire krnl_globalSort_L1_L2_11__ap_start;
  wire krnl_globalSort_L1_L2_11__ap_ready;
  wire krnl_globalSort_L1_L2_11__ap_done;
  wire krnl_globalSort_L1_L2_11__ap_idle;
  wire krnl_globalSort_L1_L2_12__ap_start;
  wire krnl_globalSort_L1_L2_12__ap_ready;
  wire krnl_globalSort_L1_L2_12__ap_done;
  wire krnl_globalSort_L1_L2_12__ap_idle;
  wire krnl_globalSort_L1_L2_13__ap_start;
  wire krnl_globalSort_L1_L2_13__ap_ready;
  wire krnl_globalSort_L1_L2_13__ap_done;
  wire krnl_globalSort_L1_L2_13__ap_idle;
  wire krnl_globalSort_L1_L2_14__ap_start;
  wire krnl_globalSort_L1_L2_14__ap_ready;
  wire krnl_globalSort_L1_L2_14__ap_done;
  wire krnl_globalSort_L1_L2_14__ap_idle;
  wire krnl_globalSort_L1_L2_15__ap_start;
  wire krnl_globalSort_L1_L2_15__ap_ready;
  wire krnl_globalSort_L1_L2_15__ap_done;
  wire krnl_globalSort_L1_L2_15__ap_idle;
  wire krnl_globalSort_L1_L2_16__ap_start;
  wire krnl_globalSort_L1_L2_16__ap_ready;
  wire krnl_globalSort_L1_L2_16__ap_done;
  wire krnl_globalSort_L1_L2_16__ap_idle;
  wire krnl_globalSort_L1_L2_17__ap_start;
  wire krnl_globalSort_L1_L2_17__ap_ready;
  wire krnl_globalSort_L1_L2_17__ap_done;
  wire krnl_globalSort_L1_L2_17__ap_idle;
  wire krnl_globalSort_L1_L2_18__ap_start;
  wire krnl_globalSort_L1_L2_18__ap_ready;
  wire krnl_globalSort_L1_L2_18__ap_done;
  wire krnl_globalSort_L1_L2_18__ap_idle;
  wire krnl_globalSort_L1_L2_19__ap_start;
  wire krnl_globalSort_L1_L2_19__ap_ready;
  wire krnl_globalSort_L1_L2_19__ap_done;
  wire krnl_globalSort_L1_L2_19__ap_idle;
  wire krnl_globalSort_L1_L2_20__ap_start;
  wire krnl_globalSort_L1_L2_20__ap_ready;
  wire krnl_globalSort_L1_L2_20__ap_done;
  wire krnl_globalSort_L1_L2_20__ap_idle;
  wire krnl_globalSort_L1_L2_21__ap_start;
  wire krnl_globalSort_L1_L2_21__ap_ready;
  wire krnl_globalSort_L1_L2_21__ap_done;
  wire krnl_globalSort_L1_L2_21__ap_idle;
  wire krnl_globalSort_L1_L2_22__ap_start;
  wire krnl_globalSort_L1_L2_22__ap_ready;
  wire krnl_globalSort_L1_L2_22__ap_done;
  wire krnl_globalSort_L1_L2_22__ap_idle;
  wire krnl_globalSort_L1_L2_23__ap_start;
  wire krnl_globalSort_L1_L2_23__ap_ready;
  wire krnl_globalSort_L1_L2_23__ap_done;
  wire krnl_globalSort_L1_L2_23__ap_idle;
  wire krnl_globalSort_L1_L2_24__ap_start;
  wire krnl_globalSort_L1_L2_24__ap_ready;
  wire krnl_globalSort_L1_L2_24__ap_done;
  wire krnl_globalSort_L1_L2_24__ap_idle;
  wire krnl_globalSort_L1_L2_25__ap_start;
  wire krnl_globalSort_L1_L2_25__ap_ready;
  wire krnl_globalSort_L1_L2_25__ap_done;
  wire krnl_globalSort_L1_L2_25__ap_idle;
  wire [63:0] krnl_globalSort_L3_0___L4_out_dist__q0;
  wire [63:0] L4_out_dist_read_addr__din;
  wire L4_out_dist_read_addr__full_n;
  wire L4_out_dist_read_addr__write;
  wire [31:0] L4_out_dist_read_data__dout;
  wire L4_out_dist_read_data__empty_n;
  wire L4_out_dist_read_data__read;
  wire [63:0] L4_out_dist_write_addr__din;
  wire L4_out_dist_write_addr__full_n;
  wire L4_out_dist_write_addr__write;
  wire [31:0] L4_out_dist_write_data__din;
  wire L4_out_dist_write_data__full_n;
  wire L4_out_dist_write_data__write;
  wire [7:0] L4_out_dist_write_resp__dout;
  wire L4_out_dist_write_resp__empty_n;
  wire L4_out_dist_write_resp__read;
  wire [63:0] krnl_globalSort_L3_0___L4_out_id__q0;
  wire [63:0] L4_out_id_read_addr__din;
  wire L4_out_id_read_addr__full_n;
  wire L4_out_id_read_addr__write;
  wire [31:0] L4_out_id_read_data__dout;
  wire L4_out_id_read_data__empty_n;
  wire L4_out_id_read_data__read;
  wire [63:0] L4_out_id_write_addr__din;
  wire L4_out_id_write_addr__full_n;
  wire L4_out_id_write_addr__write;
  wire [31:0] L4_out_id_write_data__din;
  wire L4_out_id_write_data__full_n;
  wire L4_out_id_write_data__write;
  wire [7:0] L4_out_id_write_resp__dout;
  wire L4_out_id_write_resp__empty_n;
  wire L4_out_id_write_resp__read;
  wire krnl_globalSort_L3_0__ap_start;
  wire krnl_globalSort_L3_0__ap_ready;
  wire krnl_globalSort_L3_0__ap_done;
  wire krnl_globalSort_L3_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_0_0___in_0__q0;
  wire [63:0] in_0_read_addr__din;
  wire in_0_read_addr__full_n;
  wire in_0_read_addr__write;
  wire [255:0] in_0_read_data__dout;
  wire in_0_read_data__empty_n;
  wire in_0_read_data__read;
  wire [63:0] in_0_write_addr__din;
  wire in_0_write_addr__full_n;
  wire in_0_write_addr__write;
  wire [255:0] in_0_write_data__din;
  wire in_0_write_data__full_n;
  wire in_0_write_data__write;
  wire [7:0] in_0_write_resp__dout;
  wire in_0_write_resp__empty_n;
  wire in_0_write_resp__read;
  wire krnl_partialKnn_wrapper_0_0__ap_start;
  wire krnl_partialKnn_wrapper_0_0__ap_ready;
  wire krnl_partialKnn_wrapper_0_0__ap_done;
  wire krnl_partialKnn_wrapper_0_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_1_0___in_1__q0;
  wire [63:0] in_1_read_addr__din;
  wire in_1_read_addr__full_n;
  wire in_1_read_addr__write;
  wire [255:0] in_1_read_data__dout;
  wire in_1_read_data__empty_n;
  wire in_1_read_data__read;
  wire [63:0] in_1_write_addr__din;
  wire in_1_write_addr__full_n;
  wire in_1_write_addr__write;
  wire [255:0] in_1_write_data__din;
  wire in_1_write_data__full_n;
  wire in_1_write_data__write;
  wire [7:0] in_1_write_resp__dout;
  wire in_1_write_resp__empty_n;
  wire in_1_write_resp__read;
  wire krnl_partialKnn_wrapper_1_0__ap_start;
  wire krnl_partialKnn_wrapper_1_0__ap_ready;
  wire krnl_partialKnn_wrapper_1_0__ap_done;
  wire krnl_partialKnn_wrapper_1_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_10_0___in_10__q0;
  wire [63:0] in_10_read_addr__din;
  wire in_10_read_addr__full_n;
  wire in_10_read_addr__write;
  wire [255:0] in_10_read_data__dout;
  wire in_10_read_data__empty_n;
  wire in_10_read_data__read;
  wire [63:0] in_10_write_addr__din;
  wire in_10_write_addr__full_n;
  wire in_10_write_addr__write;
  wire [255:0] in_10_write_data__din;
  wire in_10_write_data__full_n;
  wire in_10_write_data__write;
  wire [7:0] in_10_write_resp__dout;
  wire in_10_write_resp__empty_n;
  wire in_10_write_resp__read;
  wire krnl_partialKnn_wrapper_10_0__ap_start;
  wire krnl_partialKnn_wrapper_10_0__ap_ready;
  wire krnl_partialKnn_wrapper_10_0__ap_done;
  wire krnl_partialKnn_wrapper_10_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_11_0___in_11__q0;
  wire [63:0] in_11_read_addr__din;
  wire in_11_read_addr__full_n;
  wire in_11_read_addr__write;
  wire [255:0] in_11_read_data__dout;
  wire in_11_read_data__empty_n;
  wire in_11_read_data__read;
  wire [63:0] in_11_write_addr__din;
  wire in_11_write_addr__full_n;
  wire in_11_write_addr__write;
  wire [255:0] in_11_write_data__din;
  wire in_11_write_data__full_n;
  wire in_11_write_data__write;
  wire [7:0] in_11_write_resp__dout;
  wire in_11_write_resp__empty_n;
  wire in_11_write_resp__read;
  wire krnl_partialKnn_wrapper_11_0__ap_start;
  wire krnl_partialKnn_wrapper_11_0__ap_ready;
  wire krnl_partialKnn_wrapper_11_0__ap_done;
  wire krnl_partialKnn_wrapper_11_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_12_0___in_12__q0;
  wire [63:0] in_12_read_addr__din;
  wire in_12_read_addr__full_n;
  wire in_12_read_addr__write;
  wire [255:0] in_12_read_data__dout;
  wire in_12_read_data__empty_n;
  wire in_12_read_data__read;
  wire [63:0] in_12_write_addr__din;
  wire in_12_write_addr__full_n;
  wire in_12_write_addr__write;
  wire [255:0] in_12_write_data__din;
  wire in_12_write_data__full_n;
  wire in_12_write_data__write;
  wire [7:0] in_12_write_resp__dout;
  wire in_12_write_resp__empty_n;
  wire in_12_write_resp__read;
  wire krnl_partialKnn_wrapper_12_0__ap_start;
  wire krnl_partialKnn_wrapper_12_0__ap_ready;
  wire krnl_partialKnn_wrapper_12_0__ap_done;
  wire krnl_partialKnn_wrapper_12_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_13_0___in_13__q0;
  wire [63:0] in_13_read_addr__din;
  wire in_13_read_addr__full_n;
  wire in_13_read_addr__write;
  wire [255:0] in_13_read_data__dout;
  wire in_13_read_data__empty_n;
  wire in_13_read_data__read;
  wire [63:0] in_13_write_addr__din;
  wire in_13_write_addr__full_n;
  wire in_13_write_addr__write;
  wire [255:0] in_13_write_data__din;
  wire in_13_write_data__full_n;
  wire in_13_write_data__write;
  wire [7:0] in_13_write_resp__dout;
  wire in_13_write_resp__empty_n;
  wire in_13_write_resp__read;
  wire krnl_partialKnn_wrapper_13_0__ap_start;
  wire krnl_partialKnn_wrapper_13_0__ap_ready;
  wire krnl_partialKnn_wrapper_13_0__ap_done;
  wire krnl_partialKnn_wrapper_13_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_14_0___in_14__q0;
  wire [63:0] in_14_read_addr__din;
  wire in_14_read_addr__full_n;
  wire in_14_read_addr__write;
  wire [255:0] in_14_read_data__dout;
  wire in_14_read_data__empty_n;
  wire in_14_read_data__read;
  wire [63:0] in_14_write_addr__din;
  wire in_14_write_addr__full_n;
  wire in_14_write_addr__write;
  wire [255:0] in_14_write_data__din;
  wire in_14_write_data__full_n;
  wire in_14_write_data__write;
  wire [7:0] in_14_write_resp__dout;
  wire in_14_write_resp__empty_n;
  wire in_14_write_resp__read;
  wire krnl_partialKnn_wrapper_14_0__ap_start;
  wire krnl_partialKnn_wrapper_14_0__ap_ready;
  wire krnl_partialKnn_wrapper_14_0__ap_done;
  wire krnl_partialKnn_wrapper_14_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_15_0___in_15__q0;
  wire [63:0] in_15_read_addr__din;
  wire in_15_read_addr__full_n;
  wire in_15_read_addr__write;
  wire [255:0] in_15_read_data__dout;
  wire in_15_read_data__empty_n;
  wire in_15_read_data__read;
  wire [63:0] in_15_write_addr__din;
  wire in_15_write_addr__full_n;
  wire in_15_write_addr__write;
  wire [255:0] in_15_write_data__din;
  wire in_15_write_data__full_n;
  wire in_15_write_data__write;
  wire [7:0] in_15_write_resp__dout;
  wire in_15_write_resp__empty_n;
  wire in_15_write_resp__read;
  wire krnl_partialKnn_wrapper_15_0__ap_start;
  wire krnl_partialKnn_wrapper_15_0__ap_ready;
  wire krnl_partialKnn_wrapper_15_0__ap_done;
  wire krnl_partialKnn_wrapper_15_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_16_0___in_16__q0;
  wire [63:0] in_16_read_addr__din;
  wire in_16_read_addr__full_n;
  wire in_16_read_addr__write;
  wire [255:0] in_16_read_data__dout;
  wire in_16_read_data__empty_n;
  wire in_16_read_data__read;
  wire [63:0] in_16_write_addr__din;
  wire in_16_write_addr__full_n;
  wire in_16_write_addr__write;
  wire [255:0] in_16_write_data__din;
  wire in_16_write_data__full_n;
  wire in_16_write_data__write;
  wire [7:0] in_16_write_resp__dout;
  wire in_16_write_resp__empty_n;
  wire in_16_write_resp__read;
  wire krnl_partialKnn_wrapper_16_0__ap_start;
  wire krnl_partialKnn_wrapper_16_0__ap_ready;
  wire krnl_partialKnn_wrapper_16_0__ap_done;
  wire krnl_partialKnn_wrapper_16_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_17_0___in_17__q0;
  wire [63:0] in_17_read_addr__din;
  wire in_17_read_addr__full_n;
  wire in_17_read_addr__write;
  wire [255:0] in_17_read_data__dout;
  wire in_17_read_data__empty_n;
  wire in_17_read_data__read;
  wire [63:0] in_17_write_addr__din;
  wire in_17_write_addr__full_n;
  wire in_17_write_addr__write;
  wire [255:0] in_17_write_data__din;
  wire in_17_write_data__full_n;
  wire in_17_write_data__write;
  wire [7:0] in_17_write_resp__dout;
  wire in_17_write_resp__empty_n;
  wire in_17_write_resp__read;
  wire krnl_partialKnn_wrapper_17_0__ap_start;
  wire krnl_partialKnn_wrapper_17_0__ap_ready;
  wire krnl_partialKnn_wrapper_17_0__ap_done;
  wire krnl_partialKnn_wrapper_17_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_18_0___in_18__q0;
  wire [63:0] in_18_read_addr__din;
  wire in_18_read_addr__full_n;
  wire in_18_read_addr__write;
  wire [255:0] in_18_read_data__dout;
  wire in_18_read_data__empty_n;
  wire in_18_read_data__read;
  wire [63:0] in_18_write_addr__din;
  wire in_18_write_addr__full_n;
  wire in_18_write_addr__write;
  wire [255:0] in_18_write_data__din;
  wire in_18_write_data__full_n;
  wire in_18_write_data__write;
  wire [7:0] in_18_write_resp__dout;
  wire in_18_write_resp__empty_n;
  wire in_18_write_resp__read;
  wire krnl_partialKnn_wrapper_18_0__ap_start;
  wire krnl_partialKnn_wrapper_18_0__ap_ready;
  wire krnl_partialKnn_wrapper_18_0__ap_done;
  wire krnl_partialKnn_wrapper_18_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_19_0___in_19__q0;
  wire [63:0] in_19_read_addr__din;
  wire in_19_read_addr__full_n;
  wire in_19_read_addr__write;
  wire [255:0] in_19_read_data__dout;
  wire in_19_read_data__empty_n;
  wire in_19_read_data__read;
  wire [63:0] in_19_write_addr__din;
  wire in_19_write_addr__full_n;
  wire in_19_write_addr__write;
  wire [255:0] in_19_write_data__din;
  wire in_19_write_data__full_n;
  wire in_19_write_data__write;
  wire [7:0] in_19_write_resp__dout;
  wire in_19_write_resp__empty_n;
  wire in_19_write_resp__read;
  wire krnl_partialKnn_wrapper_19_0__ap_start;
  wire krnl_partialKnn_wrapper_19_0__ap_ready;
  wire krnl_partialKnn_wrapper_19_0__ap_done;
  wire krnl_partialKnn_wrapper_19_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_2_0___in_2__q0;
  wire [63:0] in_2_read_addr__din;
  wire in_2_read_addr__full_n;
  wire in_2_read_addr__write;
  wire [255:0] in_2_read_data__dout;
  wire in_2_read_data__empty_n;
  wire in_2_read_data__read;
  wire [63:0] in_2_write_addr__din;
  wire in_2_write_addr__full_n;
  wire in_2_write_addr__write;
  wire [255:0] in_2_write_data__din;
  wire in_2_write_data__full_n;
  wire in_2_write_data__write;
  wire [7:0] in_2_write_resp__dout;
  wire in_2_write_resp__empty_n;
  wire in_2_write_resp__read;
  wire krnl_partialKnn_wrapper_2_0__ap_start;
  wire krnl_partialKnn_wrapper_2_0__ap_ready;
  wire krnl_partialKnn_wrapper_2_0__ap_done;
  wire krnl_partialKnn_wrapper_2_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_20_0___in_20__q0;
  wire [63:0] in_20_read_addr__din;
  wire in_20_read_addr__full_n;
  wire in_20_read_addr__write;
  wire [255:0] in_20_read_data__dout;
  wire in_20_read_data__empty_n;
  wire in_20_read_data__read;
  wire [63:0] in_20_write_addr__din;
  wire in_20_write_addr__full_n;
  wire in_20_write_addr__write;
  wire [255:0] in_20_write_data__din;
  wire in_20_write_data__full_n;
  wire in_20_write_data__write;
  wire [7:0] in_20_write_resp__dout;
  wire in_20_write_resp__empty_n;
  wire in_20_write_resp__read;
  wire krnl_partialKnn_wrapper_20_0__ap_start;
  wire krnl_partialKnn_wrapper_20_0__ap_ready;
  wire krnl_partialKnn_wrapper_20_0__ap_done;
  wire krnl_partialKnn_wrapper_20_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_21_0___in_21__q0;
  wire [63:0] in_21_read_addr__din;
  wire in_21_read_addr__full_n;
  wire in_21_read_addr__write;
  wire [255:0] in_21_read_data__dout;
  wire in_21_read_data__empty_n;
  wire in_21_read_data__read;
  wire [63:0] in_21_write_addr__din;
  wire in_21_write_addr__full_n;
  wire in_21_write_addr__write;
  wire [255:0] in_21_write_data__din;
  wire in_21_write_data__full_n;
  wire in_21_write_data__write;
  wire [7:0] in_21_write_resp__dout;
  wire in_21_write_resp__empty_n;
  wire in_21_write_resp__read;
  wire krnl_partialKnn_wrapper_21_0__ap_start;
  wire krnl_partialKnn_wrapper_21_0__ap_ready;
  wire krnl_partialKnn_wrapper_21_0__ap_done;
  wire krnl_partialKnn_wrapper_21_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_22_0___in_22__q0;
  wire [63:0] in_22_read_addr__din;
  wire in_22_read_addr__full_n;
  wire in_22_read_addr__write;
  wire [255:0] in_22_read_data__dout;
  wire in_22_read_data__empty_n;
  wire in_22_read_data__read;
  wire [63:0] in_22_write_addr__din;
  wire in_22_write_addr__full_n;
  wire in_22_write_addr__write;
  wire [255:0] in_22_write_data__din;
  wire in_22_write_data__full_n;
  wire in_22_write_data__write;
  wire [7:0] in_22_write_resp__dout;
  wire in_22_write_resp__empty_n;
  wire in_22_write_resp__read;
  wire krnl_partialKnn_wrapper_22_0__ap_start;
  wire krnl_partialKnn_wrapper_22_0__ap_ready;
  wire krnl_partialKnn_wrapper_22_0__ap_done;
  wire krnl_partialKnn_wrapper_22_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_23_0___in_23__q0;
  wire [63:0] in_23_read_addr__din;
  wire in_23_read_addr__full_n;
  wire in_23_read_addr__write;
  wire [255:0] in_23_read_data__dout;
  wire in_23_read_data__empty_n;
  wire in_23_read_data__read;
  wire [63:0] in_23_write_addr__din;
  wire in_23_write_addr__full_n;
  wire in_23_write_addr__write;
  wire [255:0] in_23_write_data__din;
  wire in_23_write_data__full_n;
  wire in_23_write_data__write;
  wire [7:0] in_23_write_resp__dout;
  wire in_23_write_resp__empty_n;
  wire in_23_write_resp__read;
  wire krnl_partialKnn_wrapper_23_0__ap_start;
  wire krnl_partialKnn_wrapper_23_0__ap_ready;
  wire krnl_partialKnn_wrapper_23_0__ap_done;
  wire krnl_partialKnn_wrapper_23_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_24_0___in_24__q0;
  wire [63:0] in_24_read_addr__din;
  wire in_24_read_addr__full_n;
  wire in_24_read_addr__write;
  wire [255:0] in_24_read_data__dout;
  wire in_24_read_data__empty_n;
  wire in_24_read_data__read;
  wire [63:0] in_24_write_addr__din;
  wire in_24_write_addr__full_n;
  wire in_24_write_addr__write;
  wire [255:0] in_24_write_data__din;
  wire in_24_write_data__full_n;
  wire in_24_write_data__write;
  wire [7:0] in_24_write_resp__dout;
  wire in_24_write_resp__empty_n;
  wire in_24_write_resp__read;
  wire krnl_partialKnn_wrapper_24_0__ap_start;
  wire krnl_partialKnn_wrapper_24_0__ap_ready;
  wire krnl_partialKnn_wrapper_24_0__ap_done;
  wire krnl_partialKnn_wrapper_24_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_25_0___in_25__q0;
  wire [63:0] in_25_read_addr__din;
  wire in_25_read_addr__full_n;
  wire in_25_read_addr__write;
  wire [255:0] in_25_read_data__dout;
  wire in_25_read_data__empty_n;
  wire in_25_read_data__read;
  wire [63:0] in_25_write_addr__din;
  wire in_25_write_addr__full_n;
  wire in_25_write_addr__write;
  wire [255:0] in_25_write_data__din;
  wire in_25_write_data__full_n;
  wire in_25_write_data__write;
  wire [7:0] in_25_write_resp__dout;
  wire in_25_write_resp__empty_n;
  wire in_25_write_resp__read;
  wire krnl_partialKnn_wrapper_25_0__ap_start;
  wire krnl_partialKnn_wrapper_25_0__ap_ready;
  wire krnl_partialKnn_wrapper_25_0__ap_done;
  wire krnl_partialKnn_wrapper_25_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_26_0___in_26__q0;
  wire [63:0] in_26_read_addr__din;
  wire in_26_read_addr__full_n;
  wire in_26_read_addr__write;
  wire [255:0] in_26_read_data__dout;
  wire in_26_read_data__empty_n;
  wire in_26_read_data__read;
  wire [63:0] in_26_write_addr__din;
  wire in_26_write_addr__full_n;
  wire in_26_write_addr__write;
  wire [255:0] in_26_write_data__din;
  wire in_26_write_data__full_n;
  wire in_26_write_data__write;
  wire [7:0] in_26_write_resp__dout;
  wire in_26_write_resp__empty_n;
  wire in_26_write_resp__read;
  wire krnl_partialKnn_wrapper_26_0__ap_start;
  wire krnl_partialKnn_wrapper_26_0__ap_ready;
  wire krnl_partialKnn_wrapper_26_0__ap_done;
  wire krnl_partialKnn_wrapper_26_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_27_0___in_27__q0;
  wire [63:0] in_27_read_addr__din;
  wire in_27_read_addr__full_n;
  wire in_27_read_addr__write;
  wire [255:0] in_27_read_data__dout;
  wire in_27_read_data__empty_n;
  wire in_27_read_data__read;
  wire [63:0] in_27_write_addr__din;
  wire in_27_write_addr__full_n;
  wire in_27_write_addr__write;
  wire [255:0] in_27_write_data__din;
  wire in_27_write_data__full_n;
  wire in_27_write_data__write;
  wire [7:0] in_27_write_resp__dout;
  wire in_27_write_resp__empty_n;
  wire in_27_write_resp__read;
  wire krnl_partialKnn_wrapper_27_0__ap_start;
  wire krnl_partialKnn_wrapper_27_0__ap_ready;
  wire krnl_partialKnn_wrapper_27_0__ap_done;
  wire krnl_partialKnn_wrapper_27_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_28_0___in_28__q0;
  wire [63:0] in_28_read_addr__din;
  wire in_28_read_addr__full_n;
  wire in_28_read_addr__write;
  wire [255:0] in_28_read_data__dout;
  wire in_28_read_data__empty_n;
  wire in_28_read_data__read;
  wire [63:0] in_28_write_addr__din;
  wire in_28_write_addr__full_n;
  wire in_28_write_addr__write;
  wire [255:0] in_28_write_data__din;
  wire in_28_write_data__full_n;
  wire in_28_write_data__write;
  wire [7:0] in_28_write_resp__dout;
  wire in_28_write_resp__empty_n;
  wire in_28_write_resp__read;
  wire krnl_partialKnn_wrapper_28_0__ap_start;
  wire krnl_partialKnn_wrapper_28_0__ap_ready;
  wire krnl_partialKnn_wrapper_28_0__ap_done;
  wire krnl_partialKnn_wrapper_28_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_29_0___in_29__q0;
  wire [63:0] in_29_read_addr__din;
  wire in_29_read_addr__full_n;
  wire in_29_read_addr__write;
  wire [255:0] in_29_read_data__dout;
  wire in_29_read_data__empty_n;
  wire in_29_read_data__read;
  wire [63:0] in_29_write_addr__din;
  wire in_29_write_addr__full_n;
  wire in_29_write_addr__write;
  wire [255:0] in_29_write_data__din;
  wire in_29_write_data__full_n;
  wire in_29_write_data__write;
  wire [7:0] in_29_write_resp__dout;
  wire in_29_write_resp__empty_n;
  wire in_29_write_resp__read;
  wire krnl_partialKnn_wrapper_29_0__ap_start;
  wire krnl_partialKnn_wrapper_29_0__ap_ready;
  wire krnl_partialKnn_wrapper_29_0__ap_done;
  wire krnl_partialKnn_wrapper_29_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_3_0___in_3__q0;
  wire [63:0] in_3_read_addr__din;
  wire in_3_read_addr__full_n;
  wire in_3_read_addr__write;
  wire [255:0] in_3_read_data__dout;
  wire in_3_read_data__empty_n;
  wire in_3_read_data__read;
  wire [63:0] in_3_write_addr__din;
  wire in_3_write_addr__full_n;
  wire in_3_write_addr__write;
  wire [255:0] in_3_write_data__din;
  wire in_3_write_data__full_n;
  wire in_3_write_data__write;
  wire [7:0] in_3_write_resp__dout;
  wire in_3_write_resp__empty_n;
  wire in_3_write_resp__read;
  wire krnl_partialKnn_wrapper_3_0__ap_start;
  wire krnl_partialKnn_wrapper_3_0__ap_ready;
  wire krnl_partialKnn_wrapper_3_0__ap_done;
  wire krnl_partialKnn_wrapper_3_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_30_0___in_30__q0;
  wire [63:0] in_30_read_addr__din;
  wire in_30_read_addr__full_n;
  wire in_30_read_addr__write;
  wire [255:0] in_30_read_data__dout;
  wire in_30_read_data__empty_n;
  wire in_30_read_data__read;
  wire [63:0] in_30_write_addr__din;
  wire in_30_write_addr__full_n;
  wire in_30_write_addr__write;
  wire [255:0] in_30_write_data__din;
  wire in_30_write_data__full_n;
  wire in_30_write_data__write;
  wire [7:0] in_30_write_resp__dout;
  wire in_30_write_resp__empty_n;
  wire in_30_write_resp__read;
  wire krnl_partialKnn_wrapper_30_0__ap_start;
  wire krnl_partialKnn_wrapper_30_0__ap_ready;
  wire krnl_partialKnn_wrapper_30_0__ap_done;
  wire krnl_partialKnn_wrapper_30_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_31_0___in_31__q0;
  wire [63:0] in_31_read_addr__din;
  wire in_31_read_addr__full_n;
  wire in_31_read_addr__write;
  wire [255:0] in_31_read_data__dout;
  wire in_31_read_data__empty_n;
  wire in_31_read_data__read;
  wire [63:0] in_31_write_addr__din;
  wire in_31_write_addr__full_n;
  wire in_31_write_addr__write;
  wire [255:0] in_31_write_data__din;
  wire in_31_write_data__full_n;
  wire in_31_write_data__write;
  wire [7:0] in_31_write_resp__dout;
  wire in_31_write_resp__empty_n;
  wire in_31_write_resp__read;
  wire krnl_partialKnn_wrapper_31_0__ap_start;
  wire krnl_partialKnn_wrapper_31_0__ap_ready;
  wire krnl_partialKnn_wrapper_31_0__ap_done;
  wire krnl_partialKnn_wrapper_31_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_32_0___in_32__q0;
  wire [63:0] in_32_read_addr__din;
  wire in_32_read_addr__full_n;
  wire in_32_read_addr__write;
  wire [255:0] in_32_read_data__dout;
  wire in_32_read_data__empty_n;
  wire in_32_read_data__read;
  wire [63:0] in_32_write_addr__din;
  wire in_32_write_addr__full_n;
  wire in_32_write_addr__write;
  wire [255:0] in_32_write_data__din;
  wire in_32_write_data__full_n;
  wire in_32_write_data__write;
  wire [7:0] in_32_write_resp__dout;
  wire in_32_write_resp__empty_n;
  wire in_32_write_resp__read;
  wire krnl_partialKnn_wrapper_32_0__ap_start;
  wire krnl_partialKnn_wrapper_32_0__ap_ready;
  wire krnl_partialKnn_wrapper_32_0__ap_done;
  wire krnl_partialKnn_wrapper_32_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_33_0___in_33__q0;
  wire [63:0] in_33_read_addr__din;
  wire in_33_read_addr__full_n;
  wire in_33_read_addr__write;
  wire [255:0] in_33_read_data__dout;
  wire in_33_read_data__empty_n;
  wire in_33_read_data__read;
  wire [63:0] in_33_write_addr__din;
  wire in_33_write_addr__full_n;
  wire in_33_write_addr__write;
  wire [255:0] in_33_write_data__din;
  wire in_33_write_data__full_n;
  wire in_33_write_data__write;
  wire [7:0] in_33_write_resp__dout;
  wire in_33_write_resp__empty_n;
  wire in_33_write_resp__read;
  wire krnl_partialKnn_wrapper_33_0__ap_start;
  wire krnl_partialKnn_wrapper_33_0__ap_ready;
  wire krnl_partialKnn_wrapper_33_0__ap_done;
  wire krnl_partialKnn_wrapper_33_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_34_0___in_34__q0;
  wire [63:0] in_34_read_addr__din;
  wire in_34_read_addr__full_n;
  wire in_34_read_addr__write;
  wire [255:0] in_34_read_data__dout;
  wire in_34_read_data__empty_n;
  wire in_34_read_data__read;
  wire [63:0] in_34_write_addr__din;
  wire in_34_write_addr__full_n;
  wire in_34_write_addr__write;
  wire [255:0] in_34_write_data__din;
  wire in_34_write_data__full_n;
  wire in_34_write_data__write;
  wire [7:0] in_34_write_resp__dout;
  wire in_34_write_resp__empty_n;
  wire in_34_write_resp__read;
  wire krnl_partialKnn_wrapper_34_0__ap_start;
  wire krnl_partialKnn_wrapper_34_0__ap_ready;
  wire krnl_partialKnn_wrapper_34_0__ap_done;
  wire krnl_partialKnn_wrapper_34_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_35_0___in_35__q0;
  wire [63:0] in_35_read_addr__din;
  wire in_35_read_addr__full_n;
  wire in_35_read_addr__write;
  wire [255:0] in_35_read_data__dout;
  wire in_35_read_data__empty_n;
  wire in_35_read_data__read;
  wire [63:0] in_35_write_addr__din;
  wire in_35_write_addr__full_n;
  wire in_35_write_addr__write;
  wire [255:0] in_35_write_data__din;
  wire in_35_write_data__full_n;
  wire in_35_write_data__write;
  wire [7:0] in_35_write_resp__dout;
  wire in_35_write_resp__empty_n;
  wire in_35_write_resp__read;
  wire krnl_partialKnn_wrapper_35_0__ap_start;
  wire krnl_partialKnn_wrapper_35_0__ap_ready;
  wire krnl_partialKnn_wrapper_35_0__ap_done;
  wire krnl_partialKnn_wrapper_35_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_36_0___in_36__q0;
  wire [63:0] in_36_read_addr__din;
  wire in_36_read_addr__full_n;
  wire in_36_read_addr__write;
  wire [255:0] in_36_read_data__dout;
  wire in_36_read_data__empty_n;
  wire in_36_read_data__read;
  wire [63:0] in_36_write_addr__din;
  wire in_36_write_addr__full_n;
  wire in_36_write_addr__write;
  wire [255:0] in_36_write_data__din;
  wire in_36_write_data__full_n;
  wire in_36_write_data__write;
  wire [7:0] in_36_write_resp__dout;
  wire in_36_write_resp__empty_n;
  wire in_36_write_resp__read;
  wire krnl_partialKnn_wrapper_36_0__ap_start;
  wire krnl_partialKnn_wrapper_36_0__ap_ready;
  wire krnl_partialKnn_wrapper_36_0__ap_done;
  wire krnl_partialKnn_wrapper_36_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_37_0___in_37__q0;
  wire [63:0] in_37_read_addr__din;
  wire in_37_read_addr__full_n;
  wire in_37_read_addr__write;
  wire [255:0] in_37_read_data__dout;
  wire in_37_read_data__empty_n;
  wire in_37_read_data__read;
  wire [63:0] in_37_write_addr__din;
  wire in_37_write_addr__full_n;
  wire in_37_write_addr__write;
  wire [255:0] in_37_write_data__din;
  wire in_37_write_data__full_n;
  wire in_37_write_data__write;
  wire [7:0] in_37_write_resp__dout;
  wire in_37_write_resp__empty_n;
  wire in_37_write_resp__read;
  wire krnl_partialKnn_wrapper_37_0__ap_start;
  wire krnl_partialKnn_wrapper_37_0__ap_ready;
  wire krnl_partialKnn_wrapper_37_0__ap_done;
  wire krnl_partialKnn_wrapper_37_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_38_0___in_38__q0;
  wire [63:0] in_38_read_addr__din;
  wire in_38_read_addr__full_n;
  wire in_38_read_addr__write;
  wire [255:0] in_38_read_data__dout;
  wire in_38_read_data__empty_n;
  wire in_38_read_data__read;
  wire [63:0] in_38_write_addr__din;
  wire in_38_write_addr__full_n;
  wire in_38_write_addr__write;
  wire [255:0] in_38_write_data__din;
  wire in_38_write_data__full_n;
  wire in_38_write_data__write;
  wire [7:0] in_38_write_resp__dout;
  wire in_38_write_resp__empty_n;
  wire in_38_write_resp__read;
  wire krnl_partialKnn_wrapper_38_0__ap_start;
  wire krnl_partialKnn_wrapper_38_0__ap_ready;
  wire krnl_partialKnn_wrapper_38_0__ap_done;
  wire krnl_partialKnn_wrapper_38_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_39_0___in_39__q0;
  wire [63:0] in_39_read_addr__din;
  wire in_39_read_addr__full_n;
  wire in_39_read_addr__write;
  wire [255:0] in_39_read_data__dout;
  wire in_39_read_data__empty_n;
  wire in_39_read_data__read;
  wire [63:0] in_39_write_addr__din;
  wire in_39_write_addr__full_n;
  wire in_39_write_addr__write;
  wire [255:0] in_39_write_data__din;
  wire in_39_write_data__full_n;
  wire in_39_write_data__write;
  wire [7:0] in_39_write_resp__dout;
  wire in_39_write_resp__empty_n;
  wire in_39_write_resp__read;
  wire krnl_partialKnn_wrapper_39_0__ap_start;
  wire krnl_partialKnn_wrapper_39_0__ap_ready;
  wire krnl_partialKnn_wrapper_39_0__ap_done;
  wire krnl_partialKnn_wrapper_39_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_4_0___in_4__q0;
  wire [63:0] in_4_read_addr__din;
  wire in_4_read_addr__full_n;
  wire in_4_read_addr__write;
  wire [255:0] in_4_read_data__dout;
  wire in_4_read_data__empty_n;
  wire in_4_read_data__read;
  wire [63:0] in_4_write_addr__din;
  wire in_4_write_addr__full_n;
  wire in_4_write_addr__write;
  wire [255:0] in_4_write_data__din;
  wire in_4_write_data__full_n;
  wire in_4_write_data__write;
  wire [7:0] in_4_write_resp__dout;
  wire in_4_write_resp__empty_n;
  wire in_4_write_resp__read;
  wire krnl_partialKnn_wrapper_4_0__ap_start;
  wire krnl_partialKnn_wrapper_4_0__ap_ready;
  wire krnl_partialKnn_wrapper_4_0__ap_done;
  wire krnl_partialKnn_wrapper_4_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_40_0___in_40__q0;
  wire [63:0] in_40_read_addr__din;
  wire in_40_read_addr__full_n;
  wire in_40_read_addr__write;
  wire [255:0] in_40_read_data__dout;
  wire in_40_read_data__empty_n;
  wire in_40_read_data__read;
  wire [63:0] in_40_write_addr__din;
  wire in_40_write_addr__full_n;
  wire in_40_write_addr__write;
  wire [255:0] in_40_write_data__din;
  wire in_40_write_data__full_n;
  wire in_40_write_data__write;
  wire [7:0] in_40_write_resp__dout;
  wire in_40_write_resp__empty_n;
  wire in_40_write_resp__read;
  wire krnl_partialKnn_wrapper_40_0__ap_start;
  wire krnl_partialKnn_wrapper_40_0__ap_ready;
  wire krnl_partialKnn_wrapper_40_0__ap_done;
  wire krnl_partialKnn_wrapper_40_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_41_0___in_41__q0;
  wire [63:0] in_41_read_addr__din;
  wire in_41_read_addr__full_n;
  wire in_41_read_addr__write;
  wire [255:0] in_41_read_data__dout;
  wire in_41_read_data__empty_n;
  wire in_41_read_data__read;
  wire [63:0] in_41_write_addr__din;
  wire in_41_write_addr__full_n;
  wire in_41_write_addr__write;
  wire [255:0] in_41_write_data__din;
  wire in_41_write_data__full_n;
  wire in_41_write_data__write;
  wire [7:0] in_41_write_resp__dout;
  wire in_41_write_resp__empty_n;
  wire in_41_write_resp__read;
  wire krnl_partialKnn_wrapper_41_0__ap_start;
  wire krnl_partialKnn_wrapper_41_0__ap_ready;
  wire krnl_partialKnn_wrapper_41_0__ap_done;
  wire krnl_partialKnn_wrapper_41_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_42_0___in_42__q0;
  wire [63:0] in_42_read_addr__din;
  wire in_42_read_addr__full_n;
  wire in_42_read_addr__write;
  wire [255:0] in_42_read_data__dout;
  wire in_42_read_data__empty_n;
  wire in_42_read_data__read;
  wire [63:0] in_42_write_addr__din;
  wire in_42_write_addr__full_n;
  wire in_42_write_addr__write;
  wire [255:0] in_42_write_data__din;
  wire in_42_write_data__full_n;
  wire in_42_write_data__write;
  wire [7:0] in_42_write_resp__dout;
  wire in_42_write_resp__empty_n;
  wire in_42_write_resp__read;
  wire krnl_partialKnn_wrapper_42_0__ap_start;
  wire krnl_partialKnn_wrapper_42_0__ap_ready;
  wire krnl_partialKnn_wrapper_42_0__ap_done;
  wire krnl_partialKnn_wrapper_42_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_43_0___in_43__q0;
  wire [63:0] in_43_read_addr__din;
  wire in_43_read_addr__full_n;
  wire in_43_read_addr__write;
  wire [255:0] in_43_read_data__dout;
  wire in_43_read_data__empty_n;
  wire in_43_read_data__read;
  wire [63:0] in_43_write_addr__din;
  wire in_43_write_addr__full_n;
  wire in_43_write_addr__write;
  wire [255:0] in_43_write_data__din;
  wire in_43_write_data__full_n;
  wire in_43_write_data__write;
  wire [7:0] in_43_write_resp__dout;
  wire in_43_write_resp__empty_n;
  wire in_43_write_resp__read;
  wire krnl_partialKnn_wrapper_43_0__ap_start;
  wire krnl_partialKnn_wrapper_43_0__ap_ready;
  wire krnl_partialKnn_wrapper_43_0__ap_done;
  wire krnl_partialKnn_wrapper_43_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_44_0___in_44__q0;
  wire [63:0] in_44_read_addr__din;
  wire in_44_read_addr__full_n;
  wire in_44_read_addr__write;
  wire [255:0] in_44_read_data__dout;
  wire in_44_read_data__empty_n;
  wire in_44_read_data__read;
  wire [63:0] in_44_write_addr__din;
  wire in_44_write_addr__full_n;
  wire in_44_write_addr__write;
  wire [255:0] in_44_write_data__din;
  wire in_44_write_data__full_n;
  wire in_44_write_data__write;
  wire [7:0] in_44_write_resp__dout;
  wire in_44_write_resp__empty_n;
  wire in_44_write_resp__read;
  wire krnl_partialKnn_wrapper_44_0__ap_start;
  wire krnl_partialKnn_wrapper_44_0__ap_ready;
  wire krnl_partialKnn_wrapper_44_0__ap_done;
  wire krnl_partialKnn_wrapper_44_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_45_0___in_45__q0;
  wire [63:0] in_45_read_addr__din;
  wire in_45_read_addr__full_n;
  wire in_45_read_addr__write;
  wire [255:0] in_45_read_data__dout;
  wire in_45_read_data__empty_n;
  wire in_45_read_data__read;
  wire [63:0] in_45_write_addr__din;
  wire in_45_write_addr__full_n;
  wire in_45_write_addr__write;
  wire [255:0] in_45_write_data__din;
  wire in_45_write_data__full_n;
  wire in_45_write_data__write;
  wire [7:0] in_45_write_resp__dout;
  wire in_45_write_resp__empty_n;
  wire in_45_write_resp__read;
  wire krnl_partialKnn_wrapper_45_0__ap_start;
  wire krnl_partialKnn_wrapper_45_0__ap_ready;
  wire krnl_partialKnn_wrapper_45_0__ap_done;
  wire krnl_partialKnn_wrapper_45_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_46_0___in_46__q0;
  wire [63:0] in_46_read_addr__din;
  wire in_46_read_addr__full_n;
  wire in_46_read_addr__write;
  wire [255:0] in_46_read_data__dout;
  wire in_46_read_data__empty_n;
  wire in_46_read_data__read;
  wire [63:0] in_46_write_addr__din;
  wire in_46_write_addr__full_n;
  wire in_46_write_addr__write;
  wire [255:0] in_46_write_data__din;
  wire in_46_write_data__full_n;
  wire in_46_write_data__write;
  wire [7:0] in_46_write_resp__dout;
  wire in_46_write_resp__empty_n;
  wire in_46_write_resp__read;
  wire krnl_partialKnn_wrapper_46_0__ap_start;
  wire krnl_partialKnn_wrapper_46_0__ap_ready;
  wire krnl_partialKnn_wrapper_46_0__ap_done;
  wire krnl_partialKnn_wrapper_46_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_47_0___in_47__q0;
  wire [63:0] in_47_read_addr__din;
  wire in_47_read_addr__full_n;
  wire in_47_read_addr__write;
  wire [255:0] in_47_read_data__dout;
  wire in_47_read_data__empty_n;
  wire in_47_read_data__read;
  wire [63:0] in_47_write_addr__din;
  wire in_47_write_addr__full_n;
  wire in_47_write_addr__write;
  wire [255:0] in_47_write_data__din;
  wire in_47_write_data__full_n;
  wire in_47_write_data__write;
  wire [7:0] in_47_write_resp__dout;
  wire in_47_write_resp__empty_n;
  wire in_47_write_resp__read;
  wire krnl_partialKnn_wrapper_47_0__ap_start;
  wire krnl_partialKnn_wrapper_47_0__ap_ready;
  wire krnl_partialKnn_wrapper_47_0__ap_done;
  wire krnl_partialKnn_wrapper_47_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_48_0___in_48__q0;
  wire [63:0] in_48_read_addr__din;
  wire in_48_read_addr__full_n;
  wire in_48_read_addr__write;
  wire [255:0] in_48_read_data__dout;
  wire in_48_read_data__empty_n;
  wire in_48_read_data__read;
  wire [63:0] in_48_write_addr__din;
  wire in_48_write_addr__full_n;
  wire in_48_write_addr__write;
  wire [255:0] in_48_write_data__din;
  wire in_48_write_data__full_n;
  wire in_48_write_data__write;
  wire [7:0] in_48_write_resp__dout;
  wire in_48_write_resp__empty_n;
  wire in_48_write_resp__read;
  wire krnl_partialKnn_wrapper_48_0__ap_start;
  wire krnl_partialKnn_wrapper_48_0__ap_ready;
  wire krnl_partialKnn_wrapper_48_0__ap_done;
  wire krnl_partialKnn_wrapper_48_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_49_0___in_49__q0;
  wire [63:0] in_49_read_addr__din;
  wire in_49_read_addr__full_n;
  wire in_49_read_addr__write;
  wire [255:0] in_49_read_data__dout;
  wire in_49_read_data__empty_n;
  wire in_49_read_data__read;
  wire [63:0] in_49_write_addr__din;
  wire in_49_write_addr__full_n;
  wire in_49_write_addr__write;
  wire [255:0] in_49_write_data__din;
  wire in_49_write_data__full_n;
  wire in_49_write_data__write;
  wire [7:0] in_49_write_resp__dout;
  wire in_49_write_resp__empty_n;
  wire in_49_write_resp__read;
  wire krnl_partialKnn_wrapper_49_0__ap_start;
  wire krnl_partialKnn_wrapper_49_0__ap_ready;
  wire krnl_partialKnn_wrapper_49_0__ap_done;
  wire krnl_partialKnn_wrapper_49_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_5_0___in_5__q0;
  wire [63:0] in_5_read_addr__din;
  wire in_5_read_addr__full_n;
  wire in_5_read_addr__write;
  wire [255:0] in_5_read_data__dout;
  wire in_5_read_data__empty_n;
  wire in_5_read_data__read;
  wire [63:0] in_5_write_addr__din;
  wire in_5_write_addr__full_n;
  wire in_5_write_addr__write;
  wire [255:0] in_5_write_data__din;
  wire in_5_write_data__full_n;
  wire in_5_write_data__write;
  wire [7:0] in_5_write_resp__dout;
  wire in_5_write_resp__empty_n;
  wire in_5_write_resp__read;
  wire krnl_partialKnn_wrapper_5_0__ap_start;
  wire krnl_partialKnn_wrapper_5_0__ap_ready;
  wire krnl_partialKnn_wrapper_5_0__ap_done;
  wire krnl_partialKnn_wrapper_5_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_50_0___in_50__q0;
  wire [63:0] in_50_read_addr__din;
  wire in_50_read_addr__full_n;
  wire in_50_read_addr__write;
  wire [255:0] in_50_read_data__dout;
  wire in_50_read_data__empty_n;
  wire in_50_read_data__read;
  wire [63:0] in_50_write_addr__din;
  wire in_50_write_addr__full_n;
  wire in_50_write_addr__write;
  wire [255:0] in_50_write_data__din;
  wire in_50_write_data__full_n;
  wire in_50_write_data__write;
  wire [7:0] in_50_write_resp__dout;
  wire in_50_write_resp__empty_n;
  wire in_50_write_resp__read;
  wire krnl_partialKnn_wrapper_50_0__ap_start;
  wire krnl_partialKnn_wrapper_50_0__ap_ready;
  wire krnl_partialKnn_wrapper_50_0__ap_done;
  wire krnl_partialKnn_wrapper_50_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_51_0___in_51__q0;
  wire [63:0] in_51_read_addr__din;
  wire in_51_read_addr__full_n;
  wire in_51_read_addr__write;
  wire [255:0] in_51_read_data__dout;
  wire in_51_read_data__empty_n;
  wire in_51_read_data__read;
  wire [63:0] in_51_write_addr__din;
  wire in_51_write_addr__full_n;
  wire in_51_write_addr__write;
  wire [255:0] in_51_write_data__din;
  wire in_51_write_data__full_n;
  wire in_51_write_data__write;
  wire [7:0] in_51_write_resp__dout;
  wire in_51_write_resp__empty_n;
  wire in_51_write_resp__read;
  wire krnl_partialKnn_wrapper_51_0__ap_start;
  wire krnl_partialKnn_wrapper_51_0__ap_ready;
  wire krnl_partialKnn_wrapper_51_0__ap_done;
  wire krnl_partialKnn_wrapper_51_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_52_0___in_52__q0;
  wire [63:0] in_52_read_addr__din;
  wire in_52_read_addr__full_n;
  wire in_52_read_addr__write;
  wire [255:0] in_52_read_data__dout;
  wire in_52_read_data__empty_n;
  wire in_52_read_data__read;
  wire [63:0] in_52_write_addr__din;
  wire in_52_write_addr__full_n;
  wire in_52_write_addr__write;
  wire [255:0] in_52_write_data__din;
  wire in_52_write_data__full_n;
  wire in_52_write_data__write;
  wire [7:0] in_52_write_resp__dout;
  wire in_52_write_resp__empty_n;
  wire in_52_write_resp__read;
  wire krnl_partialKnn_wrapper_52_0__ap_start;
  wire krnl_partialKnn_wrapper_52_0__ap_ready;
  wire krnl_partialKnn_wrapper_52_0__ap_done;
  wire krnl_partialKnn_wrapper_52_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_53_0___in_53__q0;
  wire [63:0] in_53_read_addr__din;
  wire in_53_read_addr__full_n;
  wire in_53_read_addr__write;
  wire [255:0] in_53_read_data__dout;
  wire in_53_read_data__empty_n;
  wire in_53_read_data__read;
  wire [63:0] in_53_write_addr__din;
  wire in_53_write_addr__full_n;
  wire in_53_write_addr__write;
  wire [255:0] in_53_write_data__din;
  wire in_53_write_data__full_n;
  wire in_53_write_data__write;
  wire [7:0] in_53_write_resp__dout;
  wire in_53_write_resp__empty_n;
  wire in_53_write_resp__read;
  wire krnl_partialKnn_wrapper_53_0__ap_start;
  wire krnl_partialKnn_wrapper_53_0__ap_ready;
  wire krnl_partialKnn_wrapper_53_0__ap_done;
  wire krnl_partialKnn_wrapper_53_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_6_0___in_6__q0;
  wire [63:0] in_6_read_addr__din;
  wire in_6_read_addr__full_n;
  wire in_6_read_addr__write;
  wire [255:0] in_6_read_data__dout;
  wire in_6_read_data__empty_n;
  wire in_6_read_data__read;
  wire [63:0] in_6_write_addr__din;
  wire in_6_write_addr__full_n;
  wire in_6_write_addr__write;
  wire [255:0] in_6_write_data__din;
  wire in_6_write_data__full_n;
  wire in_6_write_data__write;
  wire [7:0] in_6_write_resp__dout;
  wire in_6_write_resp__empty_n;
  wire in_6_write_resp__read;
  wire krnl_partialKnn_wrapper_6_0__ap_start;
  wire krnl_partialKnn_wrapper_6_0__ap_ready;
  wire krnl_partialKnn_wrapper_6_0__ap_done;
  wire krnl_partialKnn_wrapper_6_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_7_0___in_7__q0;
  wire [63:0] in_7_read_addr__din;
  wire in_7_read_addr__full_n;
  wire in_7_read_addr__write;
  wire [255:0] in_7_read_data__dout;
  wire in_7_read_data__empty_n;
  wire in_7_read_data__read;
  wire [63:0] in_7_write_addr__din;
  wire in_7_write_addr__full_n;
  wire in_7_write_addr__write;
  wire [255:0] in_7_write_data__din;
  wire in_7_write_data__full_n;
  wire in_7_write_data__write;
  wire [7:0] in_7_write_resp__dout;
  wire in_7_write_resp__empty_n;
  wire in_7_write_resp__read;
  wire krnl_partialKnn_wrapper_7_0__ap_start;
  wire krnl_partialKnn_wrapper_7_0__ap_ready;
  wire krnl_partialKnn_wrapper_7_0__ap_done;
  wire krnl_partialKnn_wrapper_7_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_8_0___in_8__q0;
  wire [63:0] in_8_read_addr__din;
  wire in_8_read_addr__full_n;
  wire in_8_read_addr__write;
  wire [255:0] in_8_read_data__dout;
  wire in_8_read_data__empty_n;
  wire in_8_read_data__read;
  wire [63:0] in_8_write_addr__din;
  wire in_8_write_addr__full_n;
  wire in_8_write_addr__write;
  wire [255:0] in_8_write_data__din;
  wire in_8_write_data__full_n;
  wire in_8_write_data__write;
  wire [7:0] in_8_write_resp__dout;
  wire in_8_write_resp__empty_n;
  wire in_8_write_resp__read;
  wire krnl_partialKnn_wrapper_8_0__ap_start;
  wire krnl_partialKnn_wrapper_8_0__ap_ready;
  wire krnl_partialKnn_wrapper_8_0__ap_done;
  wire krnl_partialKnn_wrapper_8_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_9_0___in_9__q0;
  wire [63:0] in_9_read_addr__din;
  wire in_9_read_addr__full_n;
  wire in_9_read_addr__write;
  wire [255:0] in_9_read_data__dout;
  wire in_9_read_data__empty_n;
  wire in_9_read_data__read;
  wire [63:0] in_9_write_addr__din;
  wire in_9_write_addr__full_n;
  wire in_9_write_addr__write;
  wire [255:0] in_9_write_data__din;
  wire in_9_write_data__full_n;
  wire in_9_write_data__write;
  wire [7:0] in_9_write_resp__dout;
  wire in_9_write_resp__empty_n;
  wire in_9_write_resp__read;
  wire krnl_partialKnn_wrapper_9_0__ap_start;
  wire krnl_partialKnn_wrapper_9_0__ap_ready;
  wire krnl_partialKnn_wrapper_9_0__ap_done;
  wire krnl_partialKnn_wrapper_9_0__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  Knn_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .in_0(in_0),
    .in_1(in_1),
    .in_2(in_2),
    .in_3(in_3),
    .in_4(in_4),
    .in_5(in_5),
    .in_6(in_6),
    .in_7(in_7),
    .in_8(in_8),
    .in_9(in_9),
    .in_10(in_10),
    .in_11(in_11),
    .in_12(in_12),
    .in_13(in_13),
    .in_14(in_14),
    .in_15(in_15),
    .in_16(in_16),
    .in_17(in_17),
    .in_18(in_18),
    .in_19(in_19),
    .in_20(in_20),
    .in_21(in_21),
    .in_22(in_22),
    .in_23(in_23),
    .in_24(in_24),
    .in_25(in_25),
    .in_26(in_26),
    .in_27(in_27),
    .in_28(in_28),
    .in_29(in_29),
    .in_30(in_30),
    .in_31(in_31),
    .in_32(in_32),
    .in_33(in_33),
    .in_34(in_34),
    .in_35(in_35),
    .in_36(in_36),
    .in_37(in_37),
    .in_38(in_38),
    .in_39(in_39),
    .in_40(in_40),
    .in_41(in_41),
    .in_42(in_42),
    .in_43(in_43),
    .in_44(in_44),
    .in_45(in_45),
    .in_46(in_46),
    .in_47(in_47),
    .in_48(in_48),
    .in_49(in_49),
    .in_50(in_50),
    .in_51(in_51),
    .in_52(in_52),
    .in_53(in_53),
    .L4_out_dist(L4_out_dist),
    .L4_out_id(L4_out_id),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_0__dout),
    .if_empty_n(L1_out_dist_0__empty_n),
    .if_read(L1_out_dist_0__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_0__din),
    .if_full_n(L1_out_dist_0__full_n),
    .if_write(L1_out_dist_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_10__dout),
    .if_empty_n(L1_out_dist_10__empty_n),
    .if_read(L1_out_dist_10__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_10__din),
    .if_full_n(L1_out_dist_10__full_n),
    .if_write(L1_out_dist_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_11__dout),
    .if_empty_n(L1_out_dist_11__empty_n),
    .if_read(L1_out_dist_11__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_11__din),
    .if_full_n(L1_out_dist_11__full_n),
    .if_write(L1_out_dist_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_12__dout),
    .if_empty_n(L1_out_dist_12__empty_n),
    .if_read(L1_out_dist_12__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_12__din),
    .if_full_n(L1_out_dist_12__full_n),
    .if_write(L1_out_dist_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_13__dout),
    .if_empty_n(L1_out_dist_13__empty_n),
    .if_read(L1_out_dist_13__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_13__din),
    .if_full_n(L1_out_dist_13__full_n),
    .if_write(L1_out_dist_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_14__dout),
    .if_empty_n(L1_out_dist_14__empty_n),
    .if_read(L1_out_dist_14__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_14__din),
    .if_full_n(L1_out_dist_14__full_n),
    .if_write(L1_out_dist_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_15__dout),
    .if_empty_n(L1_out_dist_15__empty_n),
    .if_read(L1_out_dist_15__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_15__din),
    .if_full_n(L1_out_dist_15__full_n),
    .if_write(L1_out_dist_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_16__dout),
    .if_empty_n(L1_out_dist_16__empty_n),
    .if_read(L1_out_dist_16__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_16__din),
    .if_full_n(L1_out_dist_16__full_n),
    .if_write(L1_out_dist_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_17__dout),
    .if_empty_n(L1_out_dist_17__empty_n),
    .if_read(L1_out_dist_17__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_17__din),
    .if_full_n(L1_out_dist_17__full_n),
    .if_write(L1_out_dist_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_1__dout),
    .if_empty_n(L1_out_dist_1__empty_n),
    .if_read(L1_out_dist_1__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_1__din),
    .if_full_n(L1_out_dist_1__full_n),
    .if_write(L1_out_dist_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_2__dout),
    .if_empty_n(L1_out_dist_2__empty_n),
    .if_read(L1_out_dist_2__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_2__din),
    .if_full_n(L1_out_dist_2__full_n),
    .if_write(L1_out_dist_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_3__dout),
    .if_empty_n(L1_out_dist_3__empty_n),
    .if_read(L1_out_dist_3__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_3__din),
    .if_full_n(L1_out_dist_3__full_n),
    .if_write(L1_out_dist_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_4__dout),
    .if_empty_n(L1_out_dist_4__empty_n),
    .if_read(L1_out_dist_4__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_4__din),
    .if_full_n(L1_out_dist_4__full_n),
    .if_write(L1_out_dist_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_5__dout),
    .if_empty_n(L1_out_dist_5__empty_n),
    .if_read(L1_out_dist_5__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_5__din),
    .if_full_n(L1_out_dist_5__full_n),
    .if_write(L1_out_dist_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_6__dout),
    .if_empty_n(L1_out_dist_6__empty_n),
    .if_read(L1_out_dist_6__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_6__din),
    .if_full_n(L1_out_dist_6__full_n),
    .if_write(L1_out_dist_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_7__dout),
    .if_empty_n(L1_out_dist_7__empty_n),
    .if_read(L1_out_dist_7__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_7__din),
    .if_full_n(L1_out_dist_7__full_n),
    .if_write(L1_out_dist_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_8__dout),
    .if_empty_n(L1_out_dist_8__empty_n),
    .if_read(L1_out_dist_8__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_8__din),
    .if_full_n(L1_out_dist_8__full_n),
    .if_write(L1_out_dist_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_9__dout),
    .if_empty_n(L1_out_dist_9__empty_n),
    .if_read(L1_out_dist_9__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_9__din),
    .if_full_n(L1_out_dist_9__full_n),
    .if_write(L1_out_dist_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_0__dout),
    .if_empty_n(L1_out_id_0__empty_n),
    .if_read(L1_out_id_0__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_0__din),
    .if_full_n(L1_out_id_0__full_n),
    .if_write(L1_out_id_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_10__dout),
    .if_empty_n(L1_out_id_10__empty_n),
    .if_read(L1_out_id_10__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_10__din),
    .if_full_n(L1_out_id_10__full_n),
    .if_write(L1_out_id_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_11__dout),
    .if_empty_n(L1_out_id_11__empty_n),
    .if_read(L1_out_id_11__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_11__din),
    .if_full_n(L1_out_id_11__full_n),
    .if_write(L1_out_id_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_12__dout),
    .if_empty_n(L1_out_id_12__empty_n),
    .if_read(L1_out_id_12__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_12__din),
    .if_full_n(L1_out_id_12__full_n),
    .if_write(L1_out_id_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_13__dout),
    .if_empty_n(L1_out_id_13__empty_n),
    .if_read(L1_out_id_13__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_13__din),
    .if_full_n(L1_out_id_13__full_n),
    .if_write(L1_out_id_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_14__dout),
    .if_empty_n(L1_out_id_14__empty_n),
    .if_read(L1_out_id_14__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_14__din),
    .if_full_n(L1_out_id_14__full_n),
    .if_write(L1_out_id_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_15__dout),
    .if_empty_n(L1_out_id_15__empty_n),
    .if_read(L1_out_id_15__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_15__din),
    .if_full_n(L1_out_id_15__full_n),
    .if_write(L1_out_id_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_16__dout),
    .if_empty_n(L1_out_id_16__empty_n),
    .if_read(L1_out_id_16__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_16__din),
    .if_full_n(L1_out_id_16__full_n),
    .if_write(L1_out_id_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_17__dout),
    .if_empty_n(L1_out_id_17__empty_n),
    .if_read(L1_out_id_17__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_17__din),
    .if_full_n(L1_out_id_17__full_n),
    .if_write(L1_out_id_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_1__dout),
    .if_empty_n(L1_out_id_1__empty_n),
    .if_read(L1_out_id_1__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_1__din),
    .if_full_n(L1_out_id_1__full_n),
    .if_write(L1_out_id_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_2__dout),
    .if_empty_n(L1_out_id_2__empty_n),
    .if_read(L1_out_id_2__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_2__din),
    .if_full_n(L1_out_id_2__full_n),
    .if_write(L1_out_id_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_3__dout),
    .if_empty_n(L1_out_id_3__empty_n),
    .if_read(L1_out_id_3__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_3__din),
    .if_full_n(L1_out_id_3__full_n),
    .if_write(L1_out_id_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_4__dout),
    .if_empty_n(L1_out_id_4__empty_n),
    .if_read(L1_out_id_4__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_4__din),
    .if_full_n(L1_out_id_4__full_n),
    .if_write(L1_out_id_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_5__dout),
    .if_empty_n(L1_out_id_5__empty_n),
    .if_read(L1_out_id_5__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_5__din),
    .if_full_n(L1_out_id_5__full_n),
    .if_write(L1_out_id_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_6__dout),
    .if_empty_n(L1_out_id_6__empty_n),
    .if_read(L1_out_id_6__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_6__din),
    .if_full_n(L1_out_id_6__full_n),
    .if_write(L1_out_id_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_7__dout),
    .if_empty_n(L1_out_id_7__empty_n),
    .if_read(L1_out_id_7__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_7__din),
    .if_full_n(L1_out_id_7__full_n),
    .if_write(L1_out_id_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_8__dout),
    .if_empty_n(L1_out_id_8__empty_n),
    .if_read(L1_out_id_8__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_8__din),
    .if_full_n(L1_out_id_8__full_n),
    .if_write(L1_out_id_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_9__dout),
    .if_empty_n(L1_out_id_9__empty_n),
    .if_read(L1_out_id_9__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_9__din),
    .if_full_n(L1_out_id_9__full_n),
    .if_write(L1_out_id_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist0__dout),
    .if_empty_n(L2_out_dist0__empty_n),
    .if_read(L2_out_dist0__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist0__din),
    .if_full_n(L2_out_dist0__full_n),
    .if_write(L2_out_dist0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist1__dout),
    .if_empty_n(L2_out_dist1__empty_n),
    .if_read(L2_out_dist1__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist1__din),
    .if_full_n(L2_out_dist1__full_n),
    .if_write(L2_out_dist1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist2__dout),
    .if_empty_n(L2_out_dist2__empty_n),
    .if_read(L2_out_dist2__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist2__din),
    .if_full_n(L2_out_dist2__full_n),
    .if_write(L2_out_dist2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist3__dout),
    .if_empty_n(L2_out_dist3__empty_n),
    .if_read(L2_out_dist3__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist3__din),
    .if_full_n(L2_out_dist3__full_n),
    .if_write(L2_out_dist3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist4__dout),
    .if_empty_n(L2_out_dist4__empty_n),
    .if_read(L2_out_dist4__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist4__din),
    .if_full_n(L2_out_dist4__full_n),
    .if_write(L2_out_dist4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist5__dout),
    .if_empty_n(L2_out_dist5__empty_n),
    .if_read(L2_out_dist5__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist5__din),
    .if_full_n(L2_out_dist5__full_n),
    .if_write(L2_out_dist5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id0__dout),
    .if_empty_n(L2_out_id0__empty_n),
    .if_read(L2_out_id0__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id0__din),
    .if_full_n(L2_out_id0__full_n),
    .if_write(L2_out_id0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id1__dout),
    .if_empty_n(L2_out_id1__empty_n),
    .if_read(L2_out_id1__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id1__din),
    .if_full_n(L2_out_id1__full_n),
    .if_write(L2_out_id1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id2__dout),
    .if_empty_n(L2_out_id2__empty_n),
    .if_read(L2_out_id2__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id2__din),
    .if_full_n(L2_out_id2__full_n),
    .if_write(L2_out_id2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id3__dout),
    .if_empty_n(L2_out_id3__empty_n),
    .if_read(L2_out_id3__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id3__din),
    .if_full_n(L2_out_id3__full_n),
    .if_write(L2_out_id3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id4__dout),
    .if_empty_n(L2_out_id4__empty_n),
    .if_read(L2_out_id4__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id4__din),
    .if_full_n(L2_out_id4__full_n),
    .if_write(L2_out_id4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id5__dout),
    .if_empty_n(L2_out_id5__empty_n),
    .if_read(L2_out_id5__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id5__din),
    .if_full_n(L2_out_id5__full_n),
    .if_write(L2_out_id5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L3_out_dist0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L3_out_dist0__dout),
    .if_empty_n(L3_out_dist0__empty_n),
    .if_read(L3_out_dist0__read),
    .if_read_ce(1'b1),
    .if_din(L3_out_dist0__din),
    .if_full_n(L3_out_dist0__full_n),
    .if_write(L3_out_dist0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L3_out_dist1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L3_out_dist1__dout),
    .if_empty_n(L3_out_dist1__empty_n),
    .if_read(L3_out_dist1__read),
    .if_read_ce(1'b1),
    .if_din(L3_out_dist1__din),
    .if_full_n(L3_out_dist1__full_n),
    .if_write(L3_out_dist1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L3_out_id0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L3_out_id0__dout),
    .if_empty_n(L3_out_id0__empty_n),
    .if_read(L3_out_id0__read),
    .if_read_ce(1'b1),
    .if_din(L3_out_id0__din),
    .if_full_n(L3_out_id0__full_n),
    .if_write(L3_out_id0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L3_out_id1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L3_out_id1__dout),
    .if_empty_n(L3_out_id1__empty_n),
    .if_read(L3_out_id1__read),
    .if_read_ce(1'b1),
    .if_din(L3_out_id1__din),
    .if_full_n(L3_out_id1__full_n),
    .if_write(L3_out_id1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_0__dout),
    .if_empty_n(out_dist_0__empty_n),
    .if_read(out_dist_0__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_0__din),
    .if_full_n(out_dist_0__full_n),
    .if_write(out_dist_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_10__dout),
    .if_empty_n(out_dist_10__empty_n),
    .if_read(out_dist_10__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_10__din),
    .if_full_n(out_dist_10__full_n),
    .if_write(out_dist_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_11__dout),
    .if_empty_n(out_dist_11__empty_n),
    .if_read(out_dist_11__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_11__din),
    .if_full_n(out_dist_11__full_n),
    .if_write(out_dist_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_12__dout),
    .if_empty_n(out_dist_12__empty_n),
    .if_read(out_dist_12__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_12__din),
    .if_full_n(out_dist_12__full_n),
    .if_write(out_dist_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_13__dout),
    .if_empty_n(out_dist_13__empty_n),
    .if_read(out_dist_13__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_13__din),
    .if_full_n(out_dist_13__full_n),
    .if_write(out_dist_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_14__dout),
    .if_empty_n(out_dist_14__empty_n),
    .if_read(out_dist_14__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_14__din),
    .if_full_n(out_dist_14__full_n),
    .if_write(out_dist_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_15__dout),
    .if_empty_n(out_dist_15__empty_n),
    .if_read(out_dist_15__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_15__din),
    .if_full_n(out_dist_15__full_n),
    .if_write(out_dist_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_16__dout),
    .if_empty_n(out_dist_16__empty_n),
    .if_read(out_dist_16__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_16__din),
    .if_full_n(out_dist_16__full_n),
    .if_write(out_dist_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_17__dout),
    .if_empty_n(out_dist_17__empty_n),
    .if_read(out_dist_17__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_17__din),
    .if_full_n(out_dist_17__full_n),
    .if_write(out_dist_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_18__dout),
    .if_empty_n(out_dist_18__empty_n),
    .if_read(out_dist_18__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_18__din),
    .if_full_n(out_dist_18__full_n),
    .if_write(out_dist_18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_19__dout),
    .if_empty_n(out_dist_19__empty_n),
    .if_read(out_dist_19__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_19__din),
    .if_full_n(out_dist_19__full_n),
    .if_write(out_dist_19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_1__dout),
    .if_empty_n(out_dist_1__empty_n),
    .if_read(out_dist_1__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_1__din),
    .if_full_n(out_dist_1__full_n),
    .if_write(out_dist_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_20__dout),
    .if_empty_n(out_dist_20__empty_n),
    .if_read(out_dist_20__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_20__din),
    .if_full_n(out_dist_20__full_n),
    .if_write(out_dist_20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_21__dout),
    .if_empty_n(out_dist_21__empty_n),
    .if_read(out_dist_21__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_21__din),
    .if_full_n(out_dist_21__full_n),
    .if_write(out_dist_21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_22__dout),
    .if_empty_n(out_dist_22__empty_n),
    .if_read(out_dist_22__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_22__din),
    .if_full_n(out_dist_22__full_n),
    .if_write(out_dist_22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_23__dout),
    .if_empty_n(out_dist_23__empty_n),
    .if_read(out_dist_23__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_23__din),
    .if_full_n(out_dist_23__full_n),
    .if_write(out_dist_23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_24__dout),
    .if_empty_n(out_dist_24__empty_n),
    .if_read(out_dist_24__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_24__din),
    .if_full_n(out_dist_24__full_n),
    .if_write(out_dist_24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_25__dout),
    .if_empty_n(out_dist_25__empty_n),
    .if_read(out_dist_25__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_25__din),
    .if_full_n(out_dist_25__full_n),
    .if_write(out_dist_25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_26__dout),
    .if_empty_n(out_dist_26__empty_n),
    .if_read(out_dist_26__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_26__din),
    .if_full_n(out_dist_26__full_n),
    .if_write(out_dist_26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_27
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_27__dout),
    .if_empty_n(out_dist_27__empty_n),
    .if_read(out_dist_27__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_27__din),
    .if_full_n(out_dist_27__full_n),
    .if_write(out_dist_27__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_28
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_28__dout),
    .if_empty_n(out_dist_28__empty_n),
    .if_read(out_dist_28__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_28__din),
    .if_full_n(out_dist_28__full_n),
    .if_write(out_dist_28__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_29
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_29__dout),
    .if_empty_n(out_dist_29__empty_n),
    .if_read(out_dist_29__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_29__din),
    .if_full_n(out_dist_29__full_n),
    .if_write(out_dist_29__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_2__dout),
    .if_empty_n(out_dist_2__empty_n),
    .if_read(out_dist_2__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_2__din),
    .if_full_n(out_dist_2__full_n),
    .if_write(out_dist_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_30
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_30__dout),
    .if_empty_n(out_dist_30__empty_n),
    .if_read(out_dist_30__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_30__din),
    .if_full_n(out_dist_30__full_n),
    .if_write(out_dist_30__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_31
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_31__dout),
    .if_empty_n(out_dist_31__empty_n),
    .if_read(out_dist_31__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_31__din),
    .if_full_n(out_dist_31__full_n),
    .if_write(out_dist_31__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_32
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_32__dout),
    .if_empty_n(out_dist_32__empty_n),
    .if_read(out_dist_32__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_32__din),
    .if_full_n(out_dist_32__full_n),
    .if_write(out_dist_32__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_33
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_33__dout),
    .if_empty_n(out_dist_33__empty_n),
    .if_read(out_dist_33__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_33__din),
    .if_full_n(out_dist_33__full_n),
    .if_write(out_dist_33__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_34
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_34__dout),
    .if_empty_n(out_dist_34__empty_n),
    .if_read(out_dist_34__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_34__din),
    .if_full_n(out_dist_34__full_n),
    .if_write(out_dist_34__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_35
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_35__dout),
    .if_empty_n(out_dist_35__empty_n),
    .if_read(out_dist_35__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_35__din),
    .if_full_n(out_dist_35__full_n),
    .if_write(out_dist_35__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_36
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_36__dout),
    .if_empty_n(out_dist_36__empty_n),
    .if_read(out_dist_36__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_36__din),
    .if_full_n(out_dist_36__full_n),
    .if_write(out_dist_36__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_37
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_37__dout),
    .if_empty_n(out_dist_37__empty_n),
    .if_read(out_dist_37__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_37__din),
    .if_full_n(out_dist_37__full_n),
    .if_write(out_dist_37__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_38
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_38__dout),
    .if_empty_n(out_dist_38__empty_n),
    .if_read(out_dist_38__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_38__din),
    .if_full_n(out_dist_38__full_n),
    .if_write(out_dist_38__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_39
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_39__dout),
    .if_empty_n(out_dist_39__empty_n),
    .if_read(out_dist_39__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_39__din),
    .if_full_n(out_dist_39__full_n),
    .if_write(out_dist_39__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_3__dout),
    .if_empty_n(out_dist_3__empty_n),
    .if_read(out_dist_3__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_3__din),
    .if_full_n(out_dist_3__full_n),
    .if_write(out_dist_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_40
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_40__dout),
    .if_empty_n(out_dist_40__empty_n),
    .if_read(out_dist_40__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_40__din),
    .if_full_n(out_dist_40__full_n),
    .if_write(out_dist_40__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_41
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_41__dout),
    .if_empty_n(out_dist_41__empty_n),
    .if_read(out_dist_41__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_41__din),
    .if_full_n(out_dist_41__full_n),
    .if_write(out_dist_41__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_42
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_42__dout),
    .if_empty_n(out_dist_42__empty_n),
    .if_read(out_dist_42__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_42__din),
    .if_full_n(out_dist_42__full_n),
    .if_write(out_dist_42__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_43
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_43__dout),
    .if_empty_n(out_dist_43__empty_n),
    .if_read(out_dist_43__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_43__din),
    .if_full_n(out_dist_43__full_n),
    .if_write(out_dist_43__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_44
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_44__dout),
    .if_empty_n(out_dist_44__empty_n),
    .if_read(out_dist_44__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_44__din),
    .if_full_n(out_dist_44__full_n),
    .if_write(out_dist_44__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_45
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_45__dout),
    .if_empty_n(out_dist_45__empty_n),
    .if_read(out_dist_45__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_45__din),
    .if_full_n(out_dist_45__full_n),
    .if_write(out_dist_45__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_46
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_46__dout),
    .if_empty_n(out_dist_46__empty_n),
    .if_read(out_dist_46__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_46__din),
    .if_full_n(out_dist_46__full_n),
    .if_write(out_dist_46__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_47
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_47__dout),
    .if_empty_n(out_dist_47__empty_n),
    .if_read(out_dist_47__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_47__din),
    .if_full_n(out_dist_47__full_n),
    .if_write(out_dist_47__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_48
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_48__dout),
    .if_empty_n(out_dist_48__empty_n),
    .if_read(out_dist_48__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_48__din),
    .if_full_n(out_dist_48__full_n),
    .if_write(out_dist_48__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_49
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_49__dout),
    .if_empty_n(out_dist_49__empty_n),
    .if_read(out_dist_49__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_49__din),
    .if_full_n(out_dist_49__full_n),
    .if_write(out_dist_49__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_4__dout),
    .if_empty_n(out_dist_4__empty_n),
    .if_read(out_dist_4__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_4__din),
    .if_full_n(out_dist_4__full_n),
    .if_write(out_dist_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_50
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_50__dout),
    .if_empty_n(out_dist_50__empty_n),
    .if_read(out_dist_50__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_50__din),
    .if_full_n(out_dist_50__full_n),
    .if_write(out_dist_50__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_51
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_51__dout),
    .if_empty_n(out_dist_51__empty_n),
    .if_read(out_dist_51__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_51__din),
    .if_full_n(out_dist_51__full_n),
    .if_write(out_dist_51__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_52
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_52__dout),
    .if_empty_n(out_dist_52__empty_n),
    .if_read(out_dist_52__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_52__din),
    .if_full_n(out_dist_52__full_n),
    .if_write(out_dist_52__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_53
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_53__dout),
    .if_empty_n(out_dist_53__empty_n),
    .if_read(out_dist_53__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_53__din),
    .if_full_n(out_dist_53__full_n),
    .if_write(out_dist_53__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_5__dout),
    .if_empty_n(out_dist_5__empty_n),
    .if_read(out_dist_5__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_5__din),
    .if_full_n(out_dist_5__full_n),
    .if_write(out_dist_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_6__dout),
    .if_empty_n(out_dist_6__empty_n),
    .if_read(out_dist_6__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_6__din),
    .if_full_n(out_dist_6__full_n),
    .if_write(out_dist_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_7__dout),
    .if_empty_n(out_dist_7__empty_n),
    .if_read(out_dist_7__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_7__din),
    .if_full_n(out_dist_7__full_n),
    .if_write(out_dist_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_8__dout),
    .if_empty_n(out_dist_8__empty_n),
    .if_read(out_dist_8__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_8__din),
    .if_full_n(out_dist_8__full_n),
    .if_write(out_dist_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_9__dout),
    .if_empty_n(out_dist_9__empty_n),
    .if_read(out_dist_9__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_9__din),
    .if_full_n(out_dist_9__full_n),
    .if_write(out_dist_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_0__dout),
    .if_empty_n(out_id_0__empty_n),
    .if_read(out_id_0__read),
    .if_read_ce(1'b1),
    .if_din(out_id_0__din),
    .if_full_n(out_id_0__full_n),
    .if_write(out_id_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_10__dout),
    .if_empty_n(out_id_10__empty_n),
    .if_read(out_id_10__read),
    .if_read_ce(1'b1),
    .if_din(out_id_10__din),
    .if_full_n(out_id_10__full_n),
    .if_write(out_id_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_11__dout),
    .if_empty_n(out_id_11__empty_n),
    .if_read(out_id_11__read),
    .if_read_ce(1'b1),
    .if_din(out_id_11__din),
    .if_full_n(out_id_11__full_n),
    .if_write(out_id_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_12__dout),
    .if_empty_n(out_id_12__empty_n),
    .if_read(out_id_12__read),
    .if_read_ce(1'b1),
    .if_din(out_id_12__din),
    .if_full_n(out_id_12__full_n),
    .if_write(out_id_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_13__dout),
    .if_empty_n(out_id_13__empty_n),
    .if_read(out_id_13__read),
    .if_read_ce(1'b1),
    .if_din(out_id_13__din),
    .if_full_n(out_id_13__full_n),
    .if_write(out_id_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_14__dout),
    .if_empty_n(out_id_14__empty_n),
    .if_read(out_id_14__read),
    .if_read_ce(1'b1),
    .if_din(out_id_14__din),
    .if_full_n(out_id_14__full_n),
    .if_write(out_id_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_15__dout),
    .if_empty_n(out_id_15__empty_n),
    .if_read(out_id_15__read),
    .if_read_ce(1'b1),
    .if_din(out_id_15__din),
    .if_full_n(out_id_15__full_n),
    .if_write(out_id_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_16__dout),
    .if_empty_n(out_id_16__empty_n),
    .if_read(out_id_16__read),
    .if_read_ce(1'b1),
    .if_din(out_id_16__din),
    .if_full_n(out_id_16__full_n),
    .if_write(out_id_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_17__dout),
    .if_empty_n(out_id_17__empty_n),
    .if_read(out_id_17__read),
    .if_read_ce(1'b1),
    .if_din(out_id_17__din),
    .if_full_n(out_id_17__full_n),
    .if_write(out_id_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_18__dout),
    .if_empty_n(out_id_18__empty_n),
    .if_read(out_id_18__read),
    .if_read_ce(1'b1),
    .if_din(out_id_18__din),
    .if_full_n(out_id_18__full_n),
    .if_write(out_id_18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_19__dout),
    .if_empty_n(out_id_19__empty_n),
    .if_read(out_id_19__read),
    .if_read_ce(1'b1),
    .if_din(out_id_19__din),
    .if_full_n(out_id_19__full_n),
    .if_write(out_id_19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_1__dout),
    .if_empty_n(out_id_1__empty_n),
    .if_read(out_id_1__read),
    .if_read_ce(1'b1),
    .if_din(out_id_1__din),
    .if_full_n(out_id_1__full_n),
    .if_write(out_id_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_20__dout),
    .if_empty_n(out_id_20__empty_n),
    .if_read(out_id_20__read),
    .if_read_ce(1'b1),
    .if_din(out_id_20__din),
    .if_full_n(out_id_20__full_n),
    .if_write(out_id_20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_21__dout),
    .if_empty_n(out_id_21__empty_n),
    .if_read(out_id_21__read),
    .if_read_ce(1'b1),
    .if_din(out_id_21__din),
    .if_full_n(out_id_21__full_n),
    .if_write(out_id_21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_22__dout),
    .if_empty_n(out_id_22__empty_n),
    .if_read(out_id_22__read),
    .if_read_ce(1'b1),
    .if_din(out_id_22__din),
    .if_full_n(out_id_22__full_n),
    .if_write(out_id_22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_23__dout),
    .if_empty_n(out_id_23__empty_n),
    .if_read(out_id_23__read),
    .if_read_ce(1'b1),
    .if_din(out_id_23__din),
    .if_full_n(out_id_23__full_n),
    .if_write(out_id_23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_24__dout),
    .if_empty_n(out_id_24__empty_n),
    .if_read(out_id_24__read),
    .if_read_ce(1'b1),
    .if_din(out_id_24__din),
    .if_full_n(out_id_24__full_n),
    .if_write(out_id_24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_25__dout),
    .if_empty_n(out_id_25__empty_n),
    .if_read(out_id_25__read),
    .if_read_ce(1'b1),
    .if_din(out_id_25__din),
    .if_full_n(out_id_25__full_n),
    .if_write(out_id_25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_26__dout),
    .if_empty_n(out_id_26__empty_n),
    .if_read(out_id_26__read),
    .if_read_ce(1'b1),
    .if_din(out_id_26__din),
    .if_full_n(out_id_26__full_n),
    .if_write(out_id_26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_27
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_27__dout),
    .if_empty_n(out_id_27__empty_n),
    .if_read(out_id_27__read),
    .if_read_ce(1'b1),
    .if_din(out_id_27__din),
    .if_full_n(out_id_27__full_n),
    .if_write(out_id_27__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_28
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_28__dout),
    .if_empty_n(out_id_28__empty_n),
    .if_read(out_id_28__read),
    .if_read_ce(1'b1),
    .if_din(out_id_28__din),
    .if_full_n(out_id_28__full_n),
    .if_write(out_id_28__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_29
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_29__dout),
    .if_empty_n(out_id_29__empty_n),
    .if_read(out_id_29__read),
    .if_read_ce(1'b1),
    .if_din(out_id_29__din),
    .if_full_n(out_id_29__full_n),
    .if_write(out_id_29__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_2__dout),
    .if_empty_n(out_id_2__empty_n),
    .if_read(out_id_2__read),
    .if_read_ce(1'b1),
    .if_din(out_id_2__din),
    .if_full_n(out_id_2__full_n),
    .if_write(out_id_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_30
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_30__dout),
    .if_empty_n(out_id_30__empty_n),
    .if_read(out_id_30__read),
    .if_read_ce(1'b1),
    .if_din(out_id_30__din),
    .if_full_n(out_id_30__full_n),
    .if_write(out_id_30__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_31
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_31__dout),
    .if_empty_n(out_id_31__empty_n),
    .if_read(out_id_31__read),
    .if_read_ce(1'b1),
    .if_din(out_id_31__din),
    .if_full_n(out_id_31__full_n),
    .if_write(out_id_31__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_32
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_32__dout),
    .if_empty_n(out_id_32__empty_n),
    .if_read(out_id_32__read),
    .if_read_ce(1'b1),
    .if_din(out_id_32__din),
    .if_full_n(out_id_32__full_n),
    .if_write(out_id_32__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_33
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_33__dout),
    .if_empty_n(out_id_33__empty_n),
    .if_read(out_id_33__read),
    .if_read_ce(1'b1),
    .if_din(out_id_33__din),
    .if_full_n(out_id_33__full_n),
    .if_write(out_id_33__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_34
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_34__dout),
    .if_empty_n(out_id_34__empty_n),
    .if_read(out_id_34__read),
    .if_read_ce(1'b1),
    .if_din(out_id_34__din),
    .if_full_n(out_id_34__full_n),
    .if_write(out_id_34__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_35
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_35__dout),
    .if_empty_n(out_id_35__empty_n),
    .if_read(out_id_35__read),
    .if_read_ce(1'b1),
    .if_din(out_id_35__din),
    .if_full_n(out_id_35__full_n),
    .if_write(out_id_35__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_36
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_36__dout),
    .if_empty_n(out_id_36__empty_n),
    .if_read(out_id_36__read),
    .if_read_ce(1'b1),
    .if_din(out_id_36__din),
    .if_full_n(out_id_36__full_n),
    .if_write(out_id_36__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_37
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_37__dout),
    .if_empty_n(out_id_37__empty_n),
    .if_read(out_id_37__read),
    .if_read_ce(1'b1),
    .if_din(out_id_37__din),
    .if_full_n(out_id_37__full_n),
    .if_write(out_id_37__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_38
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_38__dout),
    .if_empty_n(out_id_38__empty_n),
    .if_read(out_id_38__read),
    .if_read_ce(1'b1),
    .if_din(out_id_38__din),
    .if_full_n(out_id_38__full_n),
    .if_write(out_id_38__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_39
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_39__dout),
    .if_empty_n(out_id_39__empty_n),
    .if_read(out_id_39__read),
    .if_read_ce(1'b1),
    .if_din(out_id_39__din),
    .if_full_n(out_id_39__full_n),
    .if_write(out_id_39__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_3__dout),
    .if_empty_n(out_id_3__empty_n),
    .if_read(out_id_3__read),
    .if_read_ce(1'b1),
    .if_din(out_id_3__din),
    .if_full_n(out_id_3__full_n),
    .if_write(out_id_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_40
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_40__dout),
    .if_empty_n(out_id_40__empty_n),
    .if_read(out_id_40__read),
    .if_read_ce(1'b1),
    .if_din(out_id_40__din),
    .if_full_n(out_id_40__full_n),
    .if_write(out_id_40__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_41
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_41__dout),
    .if_empty_n(out_id_41__empty_n),
    .if_read(out_id_41__read),
    .if_read_ce(1'b1),
    .if_din(out_id_41__din),
    .if_full_n(out_id_41__full_n),
    .if_write(out_id_41__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_42
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_42__dout),
    .if_empty_n(out_id_42__empty_n),
    .if_read(out_id_42__read),
    .if_read_ce(1'b1),
    .if_din(out_id_42__din),
    .if_full_n(out_id_42__full_n),
    .if_write(out_id_42__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_43
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_43__dout),
    .if_empty_n(out_id_43__empty_n),
    .if_read(out_id_43__read),
    .if_read_ce(1'b1),
    .if_din(out_id_43__din),
    .if_full_n(out_id_43__full_n),
    .if_write(out_id_43__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_44
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_44__dout),
    .if_empty_n(out_id_44__empty_n),
    .if_read(out_id_44__read),
    .if_read_ce(1'b1),
    .if_din(out_id_44__din),
    .if_full_n(out_id_44__full_n),
    .if_write(out_id_44__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_45
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_45__dout),
    .if_empty_n(out_id_45__empty_n),
    .if_read(out_id_45__read),
    .if_read_ce(1'b1),
    .if_din(out_id_45__din),
    .if_full_n(out_id_45__full_n),
    .if_write(out_id_45__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_46
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_46__dout),
    .if_empty_n(out_id_46__empty_n),
    .if_read(out_id_46__read),
    .if_read_ce(1'b1),
    .if_din(out_id_46__din),
    .if_full_n(out_id_46__full_n),
    .if_write(out_id_46__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_47
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_47__dout),
    .if_empty_n(out_id_47__empty_n),
    .if_read(out_id_47__read),
    .if_read_ce(1'b1),
    .if_din(out_id_47__din),
    .if_full_n(out_id_47__full_n),
    .if_write(out_id_47__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_48
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_48__dout),
    .if_empty_n(out_id_48__empty_n),
    .if_read(out_id_48__read),
    .if_read_ce(1'b1),
    .if_din(out_id_48__din),
    .if_full_n(out_id_48__full_n),
    .if_write(out_id_48__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_49
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_49__dout),
    .if_empty_n(out_id_49__empty_n),
    .if_read(out_id_49__read),
    .if_read_ce(1'b1),
    .if_din(out_id_49__din),
    .if_full_n(out_id_49__full_n),
    .if_write(out_id_49__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_4__dout),
    .if_empty_n(out_id_4__empty_n),
    .if_read(out_id_4__read),
    .if_read_ce(1'b1),
    .if_din(out_id_4__din),
    .if_full_n(out_id_4__full_n),
    .if_write(out_id_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_50
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_50__dout),
    .if_empty_n(out_id_50__empty_n),
    .if_read(out_id_50__read),
    .if_read_ce(1'b1),
    .if_din(out_id_50__din),
    .if_full_n(out_id_50__full_n),
    .if_write(out_id_50__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_51
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_51__dout),
    .if_empty_n(out_id_51__empty_n),
    .if_read(out_id_51__read),
    .if_read_ce(1'b1),
    .if_din(out_id_51__din),
    .if_full_n(out_id_51__full_n),
    .if_write(out_id_51__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_52
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_52__dout),
    .if_empty_n(out_id_52__empty_n),
    .if_read(out_id_52__read),
    .if_read_ce(1'b1),
    .if_din(out_id_52__din),
    .if_full_n(out_id_52__full_n),
    .if_write(out_id_52__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_53
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_53__dout),
    .if_empty_n(out_id_53__empty_n),
    .if_read(out_id_53__read),
    .if_read_ce(1'b1),
    .if_din(out_id_53__din),
    .if_full_n(out_id_53__full_n),
    .if_write(out_id_53__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_5__dout),
    .if_empty_n(out_id_5__empty_n),
    .if_read(out_id_5__read),
    .if_read_ce(1'b1),
    .if_din(out_id_5__din),
    .if_full_n(out_id_5__full_n),
    .if_write(out_id_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_6__dout),
    .if_empty_n(out_id_6__empty_n),
    .if_read(out_id_6__read),
    .if_read_ce(1'b1),
    .if_din(out_id_6__din),
    .if_full_n(out_id_6__full_n),
    .if_write(out_id_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_7__dout),
    .if_empty_n(out_id_7__empty_n),
    .if_read(out_id_7__read),
    .if_read_ce(1'b1),
    .if_din(out_id_7__din),
    .if_full_n(out_id_7__full_n),
    .if_write(out_id_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_8__dout),
    .if_empty_n(out_id_8__empty_n),
    .if_read(out_id_8__read),
    .if_read_ce(1'b1),
    .if_din(out_id_8__din),
    .if_full_n(out_id_8__full_n),
    .if_write(out_id_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_9__dout),
    .if_empty_n(out_id_9__empty_n),
    .if_read(out_id_9__read),
    .if_read_ce(1'b1),
    .if_din(out_id_9__din),
    .if_full_n(out_id_9__full_n),
    .if_write(out_id_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_0__ap_start),
    .ap_done(krnl_globalSort_L1_L2_0__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_0__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_0__ap_ready),
    .out_dist_din(L1_out_dist_0__din),
    .out_dist_full_n(L1_out_dist_0__full_n),
    .out_dist_write(L1_out_dist_0__write),
    .out_id_din(L1_out_id_0__din),
    .out_id_full_n(L1_out_id_0__full_n),
    .out_id_write(L1_out_id_0__write),
    .in_dist0_s_dout(out_dist_0__dout),
    .in_dist0_peek_dout(out_dist_0__dout),
    .in_dist0_s_empty_n(out_dist_0__empty_n),
    .in_dist0_peek_empty_n(out_dist_0__empty_n),
    .in_dist0_s_read(out_dist_0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_1__dout),
    .in_dist1_peek_dout(out_dist_1__dout),
    .in_dist1_s_empty_n(out_dist_1__empty_n),
    .in_dist1_peek_empty_n(out_dist_1__empty_n),
    .in_dist1_s_read(out_dist_1__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_2__dout),
    .in_dist2_peek_dout(out_dist_2__dout),
    .in_dist2_s_empty_n(out_dist_2__empty_n),
    .in_dist2_peek_empty_n(out_dist_2__empty_n),
    .in_dist2_s_read(out_dist_2__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_0__dout),
    .in_id0_peek_dout(out_id_0__dout),
    .in_id0_s_empty_n(out_id_0__empty_n),
    .in_id0_peek_empty_n(out_id_0__empty_n),
    .in_id0_s_read(out_id_0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_1__dout),
    .in_id1_peek_dout(out_id_1__dout),
    .in_id1_s_empty_n(out_id_1__empty_n),
    .in_id1_peek_empty_n(out_id_1__empty_n),
    .in_id1_s_read(out_id_1__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_2__dout),
    .in_id2_peek_dout(out_id_2__dout),
    .in_id2_s_empty_n(out_id_2__empty_n),
    .in_id2_peek_empty_n(out_id_2__empty_n),
    .in_id2_s_read(out_id_2__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_1__ap_start),
    .ap_done(krnl_globalSort_L1_L2_1__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_1__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_1__ap_ready),
    .out_dist_din(L1_out_dist_1__din),
    .out_dist_full_n(L1_out_dist_1__full_n),
    .out_dist_write(L1_out_dist_1__write),
    .out_id_din(L1_out_id_1__din),
    .out_id_full_n(L1_out_id_1__full_n),
    .out_id_write(L1_out_id_1__write),
    .in_dist0_s_dout(out_dist_3__dout),
    .in_dist0_peek_dout(out_dist_3__dout),
    .in_dist0_s_empty_n(out_dist_3__empty_n),
    .in_dist0_peek_empty_n(out_dist_3__empty_n),
    .in_dist0_s_read(out_dist_3__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_4__dout),
    .in_dist1_peek_dout(out_dist_4__dout),
    .in_dist1_s_empty_n(out_dist_4__empty_n),
    .in_dist1_peek_empty_n(out_dist_4__empty_n),
    .in_dist1_s_read(out_dist_4__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_5__dout),
    .in_dist2_peek_dout(out_dist_5__dout),
    .in_dist2_s_empty_n(out_dist_5__empty_n),
    .in_dist2_peek_empty_n(out_dist_5__empty_n),
    .in_dist2_s_read(out_dist_5__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_3__dout),
    .in_id0_peek_dout(out_id_3__dout),
    .in_id0_s_empty_n(out_id_3__empty_n),
    .in_id0_peek_empty_n(out_id_3__empty_n),
    .in_id0_s_read(out_id_3__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_4__dout),
    .in_id1_peek_dout(out_id_4__dout),
    .in_id1_s_empty_n(out_id_4__empty_n),
    .in_id1_peek_empty_n(out_id_4__empty_n),
    .in_id1_s_read(out_id_4__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_5__dout),
    .in_id2_peek_dout(out_id_5__dout),
    .in_id2_s_empty_n(out_id_5__empty_n),
    .in_id2_peek_empty_n(out_id_5__empty_n),
    .in_id2_s_read(out_id_5__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_2__ap_start),
    .ap_done(krnl_globalSort_L1_L2_2__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_2__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_2__ap_ready),
    .out_dist_din(L1_out_dist_2__din),
    .out_dist_full_n(L1_out_dist_2__full_n),
    .out_dist_write(L1_out_dist_2__write),
    .out_id_din(L1_out_id_2__din),
    .out_id_full_n(L1_out_id_2__full_n),
    .out_id_write(L1_out_id_2__write),
    .in_dist0_s_dout(out_dist_6__dout),
    .in_dist0_peek_dout(out_dist_6__dout),
    .in_dist0_s_empty_n(out_dist_6__empty_n),
    .in_dist0_peek_empty_n(out_dist_6__empty_n),
    .in_dist0_s_read(out_dist_6__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_7__dout),
    .in_dist1_peek_dout(out_dist_7__dout),
    .in_dist1_s_empty_n(out_dist_7__empty_n),
    .in_dist1_peek_empty_n(out_dist_7__empty_n),
    .in_dist1_s_read(out_dist_7__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_8__dout),
    .in_dist2_peek_dout(out_dist_8__dout),
    .in_dist2_s_empty_n(out_dist_8__empty_n),
    .in_dist2_peek_empty_n(out_dist_8__empty_n),
    .in_dist2_s_read(out_dist_8__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_6__dout),
    .in_id0_peek_dout(out_id_6__dout),
    .in_id0_s_empty_n(out_id_6__empty_n),
    .in_id0_peek_empty_n(out_id_6__empty_n),
    .in_id0_s_read(out_id_6__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_7__dout),
    .in_id1_peek_dout(out_id_7__dout),
    .in_id1_s_empty_n(out_id_7__empty_n),
    .in_id1_peek_empty_n(out_id_7__empty_n),
    .in_id1_s_read(out_id_7__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_8__dout),
    .in_id2_peek_dout(out_id_8__dout),
    .in_id2_s_empty_n(out_id_8__empty_n),
    .in_id2_peek_empty_n(out_id_8__empty_n),
    .in_id2_s_read(out_id_8__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_3__ap_start),
    .ap_done(krnl_globalSort_L1_L2_3__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_3__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_3__ap_ready),
    .out_dist_din(L1_out_dist_3__din),
    .out_dist_full_n(L1_out_dist_3__full_n),
    .out_dist_write(L1_out_dist_3__write),
    .out_id_din(L1_out_id_3__din),
    .out_id_full_n(L1_out_id_3__full_n),
    .out_id_write(L1_out_id_3__write),
    .in_dist1_s_dout(out_dist_10__dout),
    .in_dist1_peek_dout(out_dist_10__dout),
    .in_dist1_s_empty_n(out_dist_10__empty_n),
    .in_dist1_peek_empty_n(out_dist_10__empty_n),
    .in_dist1_s_read(out_dist_10__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_11__dout),
    .in_dist2_peek_dout(out_dist_11__dout),
    .in_dist2_s_empty_n(out_dist_11__empty_n),
    .in_dist2_peek_empty_n(out_dist_11__empty_n),
    .in_dist2_s_read(out_dist_11__read),
    .in_dist2_peek_read(),
    .in_dist0_s_dout(out_dist_9__dout),
    .in_dist0_peek_dout(out_dist_9__dout),
    .in_dist0_s_empty_n(out_dist_9__empty_n),
    .in_dist0_peek_empty_n(out_dist_9__empty_n),
    .in_dist0_s_read(out_dist_9__read),
    .in_dist0_peek_read(),
    .in_id1_s_dout(out_id_10__dout),
    .in_id1_peek_dout(out_id_10__dout),
    .in_id1_s_empty_n(out_id_10__empty_n),
    .in_id1_peek_empty_n(out_id_10__empty_n),
    .in_id1_s_read(out_id_10__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_11__dout),
    .in_id2_peek_dout(out_id_11__dout),
    .in_id2_s_empty_n(out_id_11__empty_n),
    .in_id2_peek_empty_n(out_id_11__empty_n),
    .in_id2_s_read(out_id_11__read),
    .in_id2_peek_read(),
    .in_id0_s_dout(out_id_9__dout),
    .in_id0_peek_dout(out_id_9__dout),
    .in_id0_s_empty_n(out_id_9__empty_n),
    .in_id0_peek_empty_n(out_id_9__empty_n),
    .in_id0_s_read(out_id_9__read),
    .in_id0_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_4__ap_start),
    .ap_done(krnl_globalSort_L1_L2_4__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_4__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_4__ap_ready),
    .out_dist_din(L1_out_dist_4__din),
    .out_dist_full_n(L1_out_dist_4__full_n),
    .out_dist_write(L1_out_dist_4__write),
    .out_id_din(L1_out_id_4__din),
    .out_id_full_n(L1_out_id_4__full_n),
    .out_id_write(L1_out_id_4__write),
    .in_dist0_s_dout(out_dist_12__dout),
    .in_dist0_peek_dout(out_dist_12__dout),
    .in_dist0_s_empty_n(out_dist_12__empty_n),
    .in_dist0_peek_empty_n(out_dist_12__empty_n),
    .in_dist0_s_read(out_dist_12__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_13__dout),
    .in_dist1_peek_dout(out_dist_13__dout),
    .in_dist1_s_empty_n(out_dist_13__empty_n),
    .in_dist1_peek_empty_n(out_dist_13__empty_n),
    .in_dist1_s_read(out_dist_13__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_14__dout),
    .in_dist2_peek_dout(out_dist_14__dout),
    .in_dist2_s_empty_n(out_dist_14__empty_n),
    .in_dist2_peek_empty_n(out_dist_14__empty_n),
    .in_dist2_s_read(out_dist_14__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_12__dout),
    .in_id0_peek_dout(out_id_12__dout),
    .in_id0_s_empty_n(out_id_12__empty_n),
    .in_id0_peek_empty_n(out_id_12__empty_n),
    .in_id0_s_read(out_id_12__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_13__dout),
    .in_id1_peek_dout(out_id_13__dout),
    .in_id1_s_empty_n(out_id_13__empty_n),
    .in_id1_peek_empty_n(out_id_13__empty_n),
    .in_id1_s_read(out_id_13__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_14__dout),
    .in_id2_peek_dout(out_id_14__dout),
    .in_id2_s_empty_n(out_id_14__empty_n),
    .in_id2_peek_empty_n(out_id_14__empty_n),
    .in_id2_s_read(out_id_14__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_5__ap_start),
    .ap_done(krnl_globalSort_L1_L2_5__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_5__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_5__ap_ready),
    .out_dist_din(L1_out_dist_5__din),
    .out_dist_full_n(L1_out_dist_5__full_n),
    .out_dist_write(L1_out_dist_5__write),
    .out_id_din(L1_out_id_5__din),
    .out_id_full_n(L1_out_id_5__full_n),
    .out_id_write(L1_out_id_5__write),
    .in_dist0_s_dout(out_dist_15__dout),
    .in_dist0_peek_dout(out_dist_15__dout),
    .in_dist0_s_empty_n(out_dist_15__empty_n),
    .in_dist0_peek_empty_n(out_dist_15__empty_n),
    .in_dist0_s_read(out_dist_15__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_16__dout),
    .in_dist1_peek_dout(out_dist_16__dout),
    .in_dist1_s_empty_n(out_dist_16__empty_n),
    .in_dist1_peek_empty_n(out_dist_16__empty_n),
    .in_dist1_s_read(out_dist_16__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_17__dout),
    .in_dist2_peek_dout(out_dist_17__dout),
    .in_dist2_s_empty_n(out_dist_17__empty_n),
    .in_dist2_peek_empty_n(out_dist_17__empty_n),
    .in_dist2_s_read(out_dist_17__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_15__dout),
    .in_id0_peek_dout(out_id_15__dout),
    .in_id0_s_empty_n(out_id_15__empty_n),
    .in_id0_peek_empty_n(out_id_15__empty_n),
    .in_id0_s_read(out_id_15__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_16__dout),
    .in_id1_peek_dout(out_id_16__dout),
    .in_id1_s_empty_n(out_id_16__empty_n),
    .in_id1_peek_empty_n(out_id_16__empty_n),
    .in_id1_s_read(out_id_16__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_17__dout),
    .in_id2_peek_dout(out_id_17__dout),
    .in_id2_s_empty_n(out_id_17__empty_n),
    .in_id2_peek_empty_n(out_id_17__empty_n),
    .in_id2_s_read(out_id_17__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_6__ap_start),
    .ap_done(krnl_globalSort_L1_L2_6__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_6__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_6__ap_ready),
    .out_dist_din(L1_out_dist_6__din),
    .out_dist_full_n(L1_out_dist_6__full_n),
    .out_dist_write(L1_out_dist_6__write),
    .out_id_din(L1_out_id_6__din),
    .out_id_full_n(L1_out_id_6__full_n),
    .out_id_write(L1_out_id_6__write),
    .in_dist0_s_dout(out_dist_18__dout),
    .in_dist0_peek_dout(out_dist_18__dout),
    .in_dist0_s_empty_n(out_dist_18__empty_n),
    .in_dist0_peek_empty_n(out_dist_18__empty_n),
    .in_dist0_s_read(out_dist_18__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_19__dout),
    .in_dist1_peek_dout(out_dist_19__dout),
    .in_dist1_s_empty_n(out_dist_19__empty_n),
    .in_dist1_peek_empty_n(out_dist_19__empty_n),
    .in_dist1_s_read(out_dist_19__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_20__dout),
    .in_dist2_peek_dout(out_dist_20__dout),
    .in_dist2_s_empty_n(out_dist_20__empty_n),
    .in_dist2_peek_empty_n(out_dist_20__empty_n),
    .in_dist2_s_read(out_dist_20__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_18__dout),
    .in_id0_peek_dout(out_id_18__dout),
    .in_id0_s_empty_n(out_id_18__empty_n),
    .in_id0_peek_empty_n(out_id_18__empty_n),
    .in_id0_s_read(out_id_18__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_19__dout),
    .in_id1_peek_dout(out_id_19__dout),
    .in_id1_s_empty_n(out_id_19__empty_n),
    .in_id1_peek_empty_n(out_id_19__empty_n),
    .in_id1_s_read(out_id_19__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_20__dout),
    .in_id2_peek_dout(out_id_20__dout),
    .in_id2_s_empty_n(out_id_20__empty_n),
    .in_id2_peek_empty_n(out_id_20__empty_n),
    .in_id2_s_read(out_id_20__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_7__ap_start),
    .ap_done(krnl_globalSort_L1_L2_7__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_7__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_7__ap_ready),
    .out_dist_din(L1_out_dist_7__din),
    .out_dist_full_n(L1_out_dist_7__full_n),
    .out_dist_write(L1_out_dist_7__write),
    .out_id_din(L1_out_id_7__din),
    .out_id_full_n(L1_out_id_7__full_n),
    .out_id_write(L1_out_id_7__write),
    .in_dist0_s_dout(out_dist_21__dout),
    .in_dist0_peek_dout(out_dist_21__dout),
    .in_dist0_s_empty_n(out_dist_21__empty_n),
    .in_dist0_peek_empty_n(out_dist_21__empty_n),
    .in_dist0_s_read(out_dist_21__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_22__dout),
    .in_dist1_peek_dout(out_dist_22__dout),
    .in_dist1_s_empty_n(out_dist_22__empty_n),
    .in_dist1_peek_empty_n(out_dist_22__empty_n),
    .in_dist1_s_read(out_dist_22__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_23__dout),
    .in_dist2_peek_dout(out_dist_23__dout),
    .in_dist2_s_empty_n(out_dist_23__empty_n),
    .in_dist2_peek_empty_n(out_dist_23__empty_n),
    .in_dist2_s_read(out_dist_23__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_21__dout),
    .in_id0_peek_dout(out_id_21__dout),
    .in_id0_s_empty_n(out_id_21__empty_n),
    .in_id0_peek_empty_n(out_id_21__empty_n),
    .in_id0_s_read(out_id_21__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_22__dout),
    .in_id1_peek_dout(out_id_22__dout),
    .in_id1_s_empty_n(out_id_22__empty_n),
    .in_id1_peek_empty_n(out_id_22__empty_n),
    .in_id1_s_read(out_id_22__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_23__dout),
    .in_id2_peek_dout(out_id_23__dout),
    .in_id2_s_empty_n(out_id_23__empty_n),
    .in_id2_peek_empty_n(out_id_23__empty_n),
    .in_id2_s_read(out_id_23__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_8__ap_start),
    .ap_done(krnl_globalSort_L1_L2_8__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_8__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_8__ap_ready),
    .out_dist_din(L1_out_dist_8__din),
    .out_dist_full_n(L1_out_dist_8__full_n),
    .out_dist_write(L1_out_dist_8__write),
    .out_id_din(L1_out_id_8__din),
    .out_id_full_n(L1_out_id_8__full_n),
    .out_id_write(L1_out_id_8__write),
    .in_dist0_s_dout(out_dist_24__dout),
    .in_dist0_peek_dout(out_dist_24__dout),
    .in_dist0_s_empty_n(out_dist_24__empty_n),
    .in_dist0_peek_empty_n(out_dist_24__empty_n),
    .in_dist0_s_read(out_dist_24__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_25__dout),
    .in_dist1_peek_dout(out_dist_25__dout),
    .in_dist1_s_empty_n(out_dist_25__empty_n),
    .in_dist1_peek_empty_n(out_dist_25__empty_n),
    .in_dist1_s_read(out_dist_25__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_26__dout),
    .in_dist2_peek_dout(out_dist_26__dout),
    .in_dist2_s_empty_n(out_dist_26__empty_n),
    .in_dist2_peek_empty_n(out_dist_26__empty_n),
    .in_dist2_s_read(out_dist_26__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_24__dout),
    .in_id0_peek_dout(out_id_24__dout),
    .in_id0_s_empty_n(out_id_24__empty_n),
    .in_id0_peek_empty_n(out_id_24__empty_n),
    .in_id0_s_read(out_id_24__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_25__dout),
    .in_id1_peek_dout(out_id_25__dout),
    .in_id1_s_empty_n(out_id_25__empty_n),
    .in_id1_peek_empty_n(out_id_25__empty_n),
    .in_id1_s_read(out_id_25__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_26__dout),
    .in_id2_peek_dout(out_id_26__dout),
    .in_id2_s_empty_n(out_id_26__empty_n),
    .in_id2_peek_empty_n(out_id_26__empty_n),
    .in_id2_s_read(out_id_26__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_9__ap_start),
    .ap_done(krnl_globalSort_L1_L2_9__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_9__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_9__ap_ready),
    .out_dist_din(L1_out_dist_9__din),
    .out_dist_full_n(L1_out_dist_9__full_n),
    .out_dist_write(L1_out_dist_9__write),
    .out_id_din(L1_out_id_9__din),
    .out_id_full_n(L1_out_id_9__full_n),
    .out_id_write(L1_out_id_9__write),
    .in_dist0_s_dout(out_dist_27__dout),
    .in_dist0_peek_dout(out_dist_27__dout),
    .in_dist0_s_empty_n(out_dist_27__empty_n),
    .in_dist0_peek_empty_n(out_dist_27__empty_n),
    .in_dist0_s_read(out_dist_27__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_28__dout),
    .in_dist1_peek_dout(out_dist_28__dout),
    .in_dist1_s_empty_n(out_dist_28__empty_n),
    .in_dist1_peek_empty_n(out_dist_28__empty_n),
    .in_dist1_s_read(out_dist_28__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_29__dout),
    .in_dist2_peek_dout(out_dist_29__dout),
    .in_dist2_s_empty_n(out_dist_29__empty_n),
    .in_dist2_peek_empty_n(out_dist_29__empty_n),
    .in_dist2_s_read(out_dist_29__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_27__dout),
    .in_id0_peek_dout(out_id_27__dout),
    .in_id0_s_empty_n(out_id_27__empty_n),
    .in_id0_peek_empty_n(out_id_27__empty_n),
    .in_id0_s_read(out_id_27__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_28__dout),
    .in_id1_peek_dout(out_id_28__dout),
    .in_id1_s_empty_n(out_id_28__empty_n),
    .in_id1_peek_empty_n(out_id_28__empty_n),
    .in_id1_s_read(out_id_28__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_29__dout),
    .in_id2_peek_dout(out_id_29__dout),
    .in_id2_s_empty_n(out_id_29__empty_n),
    .in_id2_peek_empty_n(out_id_29__empty_n),
    .in_id2_s_read(out_id_29__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_10__ap_start),
    .ap_done(krnl_globalSort_L1_L2_10__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_10__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_10__ap_ready),
    .out_dist_din(L1_out_dist_10__din),
    .out_dist_full_n(L1_out_dist_10__full_n),
    .out_dist_write(L1_out_dist_10__write),
    .out_id_din(L1_out_id_10__din),
    .out_id_full_n(L1_out_id_10__full_n),
    .out_id_write(L1_out_id_10__write),
    .in_dist0_s_dout(out_dist_30__dout),
    .in_dist0_peek_dout(out_dist_30__dout),
    .in_dist0_s_empty_n(out_dist_30__empty_n),
    .in_dist0_peek_empty_n(out_dist_30__empty_n),
    .in_dist0_s_read(out_dist_30__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_31__dout),
    .in_dist1_peek_dout(out_dist_31__dout),
    .in_dist1_s_empty_n(out_dist_31__empty_n),
    .in_dist1_peek_empty_n(out_dist_31__empty_n),
    .in_dist1_s_read(out_dist_31__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_32__dout),
    .in_dist2_peek_dout(out_dist_32__dout),
    .in_dist2_s_empty_n(out_dist_32__empty_n),
    .in_dist2_peek_empty_n(out_dist_32__empty_n),
    .in_dist2_s_read(out_dist_32__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_30__dout),
    .in_id0_peek_dout(out_id_30__dout),
    .in_id0_s_empty_n(out_id_30__empty_n),
    .in_id0_peek_empty_n(out_id_30__empty_n),
    .in_id0_s_read(out_id_30__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_31__dout),
    .in_id1_peek_dout(out_id_31__dout),
    .in_id1_s_empty_n(out_id_31__empty_n),
    .in_id1_peek_empty_n(out_id_31__empty_n),
    .in_id1_s_read(out_id_31__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_32__dout),
    .in_id2_peek_dout(out_id_32__dout),
    .in_id2_s_empty_n(out_id_32__empty_n),
    .in_id2_peek_empty_n(out_id_32__empty_n),
    .in_id2_s_read(out_id_32__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_11__ap_start),
    .ap_done(krnl_globalSort_L1_L2_11__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_11__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_11__ap_ready),
    .out_dist_din(L1_out_dist_11__din),
    .out_dist_full_n(L1_out_dist_11__full_n),
    .out_dist_write(L1_out_dist_11__write),
    .out_id_din(L1_out_id_11__din),
    .out_id_full_n(L1_out_id_11__full_n),
    .out_id_write(L1_out_id_11__write),
    .in_dist0_s_dout(out_dist_33__dout),
    .in_dist0_peek_dout(out_dist_33__dout),
    .in_dist0_s_empty_n(out_dist_33__empty_n),
    .in_dist0_peek_empty_n(out_dist_33__empty_n),
    .in_dist0_s_read(out_dist_33__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_34__dout),
    .in_dist1_peek_dout(out_dist_34__dout),
    .in_dist1_s_empty_n(out_dist_34__empty_n),
    .in_dist1_peek_empty_n(out_dist_34__empty_n),
    .in_dist1_s_read(out_dist_34__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_35__dout),
    .in_dist2_peek_dout(out_dist_35__dout),
    .in_dist2_s_empty_n(out_dist_35__empty_n),
    .in_dist2_peek_empty_n(out_dist_35__empty_n),
    .in_dist2_s_read(out_dist_35__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_33__dout),
    .in_id0_peek_dout(out_id_33__dout),
    .in_id0_s_empty_n(out_id_33__empty_n),
    .in_id0_peek_empty_n(out_id_33__empty_n),
    .in_id0_s_read(out_id_33__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_34__dout),
    .in_id1_peek_dout(out_id_34__dout),
    .in_id1_s_empty_n(out_id_34__empty_n),
    .in_id1_peek_empty_n(out_id_34__empty_n),
    .in_id1_s_read(out_id_34__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_35__dout),
    .in_id2_peek_dout(out_id_35__dout),
    .in_id2_s_empty_n(out_id_35__empty_n),
    .in_id2_peek_empty_n(out_id_35__empty_n),
    .in_id2_s_read(out_id_35__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_12__ap_start),
    .ap_done(krnl_globalSort_L1_L2_12__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_12__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_12__ap_ready),
    .out_dist_din(L1_out_dist_12__din),
    .out_dist_full_n(L1_out_dist_12__full_n),
    .out_dist_write(L1_out_dist_12__write),
    .out_id_din(L1_out_id_12__din),
    .out_id_full_n(L1_out_id_12__full_n),
    .out_id_write(L1_out_id_12__write),
    .in_dist0_s_dout(out_dist_36__dout),
    .in_dist0_peek_dout(out_dist_36__dout),
    .in_dist0_s_empty_n(out_dist_36__empty_n),
    .in_dist0_peek_empty_n(out_dist_36__empty_n),
    .in_dist0_s_read(out_dist_36__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_37__dout),
    .in_dist1_peek_dout(out_dist_37__dout),
    .in_dist1_s_empty_n(out_dist_37__empty_n),
    .in_dist1_peek_empty_n(out_dist_37__empty_n),
    .in_dist1_s_read(out_dist_37__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_38__dout),
    .in_dist2_peek_dout(out_dist_38__dout),
    .in_dist2_s_empty_n(out_dist_38__empty_n),
    .in_dist2_peek_empty_n(out_dist_38__empty_n),
    .in_dist2_s_read(out_dist_38__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_36__dout),
    .in_id0_peek_dout(out_id_36__dout),
    .in_id0_s_empty_n(out_id_36__empty_n),
    .in_id0_peek_empty_n(out_id_36__empty_n),
    .in_id0_s_read(out_id_36__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_37__dout),
    .in_id1_peek_dout(out_id_37__dout),
    .in_id1_s_empty_n(out_id_37__empty_n),
    .in_id1_peek_empty_n(out_id_37__empty_n),
    .in_id1_s_read(out_id_37__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_38__dout),
    .in_id2_peek_dout(out_id_38__dout),
    .in_id2_s_empty_n(out_id_38__empty_n),
    .in_id2_peek_empty_n(out_id_38__empty_n),
    .in_id2_s_read(out_id_38__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_13__ap_start),
    .ap_done(krnl_globalSort_L1_L2_13__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_13__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_13__ap_ready),
    .out_dist_din(L1_out_dist_13__din),
    .out_dist_full_n(L1_out_dist_13__full_n),
    .out_dist_write(L1_out_dist_13__write),
    .out_id_din(L1_out_id_13__din),
    .out_id_full_n(L1_out_id_13__full_n),
    .out_id_write(L1_out_id_13__write),
    .in_dist0_s_dout(out_dist_39__dout),
    .in_dist0_peek_dout(out_dist_39__dout),
    .in_dist0_s_empty_n(out_dist_39__empty_n),
    .in_dist0_peek_empty_n(out_dist_39__empty_n),
    .in_dist0_s_read(out_dist_39__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_40__dout),
    .in_dist1_peek_dout(out_dist_40__dout),
    .in_dist1_s_empty_n(out_dist_40__empty_n),
    .in_dist1_peek_empty_n(out_dist_40__empty_n),
    .in_dist1_s_read(out_dist_40__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_41__dout),
    .in_dist2_peek_dout(out_dist_41__dout),
    .in_dist2_s_empty_n(out_dist_41__empty_n),
    .in_dist2_peek_empty_n(out_dist_41__empty_n),
    .in_dist2_s_read(out_dist_41__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_39__dout),
    .in_id0_peek_dout(out_id_39__dout),
    .in_id0_s_empty_n(out_id_39__empty_n),
    .in_id0_peek_empty_n(out_id_39__empty_n),
    .in_id0_s_read(out_id_39__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_40__dout),
    .in_id1_peek_dout(out_id_40__dout),
    .in_id1_s_empty_n(out_id_40__empty_n),
    .in_id1_peek_empty_n(out_id_40__empty_n),
    .in_id1_s_read(out_id_40__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_41__dout),
    .in_id2_peek_dout(out_id_41__dout),
    .in_id2_s_empty_n(out_id_41__empty_n),
    .in_id2_peek_empty_n(out_id_41__empty_n),
    .in_id2_s_read(out_id_41__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_14__ap_start),
    .ap_done(krnl_globalSort_L1_L2_14__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_14__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_14__ap_ready),
    .out_dist_din(L1_out_dist_14__din),
    .out_dist_full_n(L1_out_dist_14__full_n),
    .out_dist_write(L1_out_dist_14__write),
    .out_id_din(L1_out_id_14__din),
    .out_id_full_n(L1_out_id_14__full_n),
    .out_id_write(L1_out_id_14__write),
    .in_dist0_s_dout(out_dist_42__dout),
    .in_dist0_peek_dout(out_dist_42__dout),
    .in_dist0_s_empty_n(out_dist_42__empty_n),
    .in_dist0_peek_empty_n(out_dist_42__empty_n),
    .in_dist0_s_read(out_dist_42__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_43__dout),
    .in_dist1_peek_dout(out_dist_43__dout),
    .in_dist1_s_empty_n(out_dist_43__empty_n),
    .in_dist1_peek_empty_n(out_dist_43__empty_n),
    .in_dist1_s_read(out_dist_43__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_44__dout),
    .in_dist2_peek_dout(out_dist_44__dout),
    .in_dist2_s_empty_n(out_dist_44__empty_n),
    .in_dist2_peek_empty_n(out_dist_44__empty_n),
    .in_dist2_s_read(out_dist_44__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_42__dout),
    .in_id0_peek_dout(out_id_42__dout),
    .in_id0_s_empty_n(out_id_42__empty_n),
    .in_id0_peek_empty_n(out_id_42__empty_n),
    .in_id0_s_read(out_id_42__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_43__dout),
    .in_id1_peek_dout(out_id_43__dout),
    .in_id1_s_empty_n(out_id_43__empty_n),
    .in_id1_peek_empty_n(out_id_43__empty_n),
    .in_id1_s_read(out_id_43__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_44__dout),
    .in_id2_peek_dout(out_id_44__dout),
    .in_id2_s_empty_n(out_id_44__empty_n),
    .in_id2_peek_empty_n(out_id_44__empty_n),
    .in_id2_s_read(out_id_44__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_15__ap_start),
    .ap_done(krnl_globalSort_L1_L2_15__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_15__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_15__ap_ready),
    .out_dist_din(L1_out_dist_15__din),
    .out_dist_full_n(L1_out_dist_15__full_n),
    .out_dist_write(L1_out_dist_15__write),
    .out_id_din(L1_out_id_15__din),
    .out_id_full_n(L1_out_id_15__full_n),
    .out_id_write(L1_out_id_15__write),
    .in_dist0_s_dout(out_dist_45__dout),
    .in_dist0_peek_dout(out_dist_45__dout),
    .in_dist0_s_empty_n(out_dist_45__empty_n),
    .in_dist0_peek_empty_n(out_dist_45__empty_n),
    .in_dist0_s_read(out_dist_45__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_46__dout),
    .in_dist1_peek_dout(out_dist_46__dout),
    .in_dist1_s_empty_n(out_dist_46__empty_n),
    .in_dist1_peek_empty_n(out_dist_46__empty_n),
    .in_dist1_s_read(out_dist_46__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_47__dout),
    .in_dist2_peek_dout(out_dist_47__dout),
    .in_dist2_s_empty_n(out_dist_47__empty_n),
    .in_dist2_peek_empty_n(out_dist_47__empty_n),
    .in_dist2_s_read(out_dist_47__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_45__dout),
    .in_id0_peek_dout(out_id_45__dout),
    .in_id0_s_empty_n(out_id_45__empty_n),
    .in_id0_peek_empty_n(out_id_45__empty_n),
    .in_id0_s_read(out_id_45__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_46__dout),
    .in_id1_peek_dout(out_id_46__dout),
    .in_id1_s_empty_n(out_id_46__empty_n),
    .in_id1_peek_empty_n(out_id_46__empty_n),
    .in_id1_s_read(out_id_46__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_47__dout),
    .in_id2_peek_dout(out_id_47__dout),
    .in_id2_s_empty_n(out_id_47__empty_n),
    .in_id2_peek_empty_n(out_id_47__empty_n),
    .in_id2_s_read(out_id_47__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_16__ap_start),
    .ap_done(krnl_globalSort_L1_L2_16__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_16__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_16__ap_ready),
    .out_dist_din(L1_out_dist_16__din),
    .out_dist_full_n(L1_out_dist_16__full_n),
    .out_dist_write(L1_out_dist_16__write),
    .out_id_din(L1_out_id_16__din),
    .out_id_full_n(L1_out_id_16__full_n),
    .out_id_write(L1_out_id_16__write),
    .in_dist0_s_dout(out_dist_48__dout),
    .in_dist0_peek_dout(out_dist_48__dout),
    .in_dist0_s_empty_n(out_dist_48__empty_n),
    .in_dist0_peek_empty_n(out_dist_48__empty_n),
    .in_dist0_s_read(out_dist_48__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_49__dout),
    .in_dist1_peek_dout(out_dist_49__dout),
    .in_dist1_s_empty_n(out_dist_49__empty_n),
    .in_dist1_peek_empty_n(out_dist_49__empty_n),
    .in_dist1_s_read(out_dist_49__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_50__dout),
    .in_dist2_peek_dout(out_dist_50__dout),
    .in_dist2_s_empty_n(out_dist_50__empty_n),
    .in_dist2_peek_empty_n(out_dist_50__empty_n),
    .in_dist2_s_read(out_dist_50__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_48__dout),
    .in_id0_peek_dout(out_id_48__dout),
    .in_id0_s_empty_n(out_id_48__empty_n),
    .in_id0_peek_empty_n(out_id_48__empty_n),
    .in_id0_s_read(out_id_48__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_49__dout),
    .in_id1_peek_dout(out_id_49__dout),
    .in_id1_s_empty_n(out_id_49__empty_n),
    .in_id1_peek_empty_n(out_id_49__empty_n),
    .in_id1_s_read(out_id_49__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_50__dout),
    .in_id2_peek_dout(out_id_50__dout),
    .in_id2_s_empty_n(out_id_50__empty_n),
    .in_id2_peek_empty_n(out_id_50__empty_n),
    .in_id2_s_read(out_id_50__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_17__ap_start),
    .ap_done(krnl_globalSort_L1_L2_17__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_17__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_17__ap_ready),
    .out_dist_din(L1_out_dist_17__din),
    .out_dist_full_n(L1_out_dist_17__full_n),
    .out_dist_write(L1_out_dist_17__write),
    .out_id_din(L1_out_id_17__din),
    .out_id_full_n(L1_out_id_17__full_n),
    .out_id_write(L1_out_id_17__write),
    .in_dist0_s_dout(out_dist_51__dout),
    .in_dist0_peek_dout(out_dist_51__dout),
    .in_dist0_s_empty_n(out_dist_51__empty_n),
    .in_dist0_peek_empty_n(out_dist_51__empty_n),
    .in_dist0_s_read(out_dist_51__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_52__dout),
    .in_dist1_peek_dout(out_dist_52__dout),
    .in_dist1_s_empty_n(out_dist_52__empty_n),
    .in_dist1_peek_empty_n(out_dist_52__empty_n),
    .in_dist1_s_read(out_dist_52__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_53__dout),
    .in_dist2_peek_dout(out_dist_53__dout),
    .in_dist2_s_empty_n(out_dist_53__empty_n),
    .in_dist2_peek_empty_n(out_dist_53__empty_n),
    .in_dist2_s_read(out_dist_53__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_51__dout),
    .in_id0_peek_dout(out_id_51__dout),
    .in_id0_s_empty_n(out_id_51__empty_n),
    .in_id0_peek_empty_n(out_id_51__empty_n),
    .in_id0_s_read(out_id_51__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_52__dout),
    .in_id1_peek_dout(out_id_52__dout),
    .in_id1_s_empty_n(out_id_52__empty_n),
    .in_id1_peek_empty_n(out_id_52__empty_n),
    .in_id1_s_read(out_id_52__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_53__dout),
    .in_id2_peek_dout(out_id_53__dout),
    .in_id2_s_empty_n(out_id_53__empty_n),
    .in_id2_peek_empty_n(out_id_53__empty_n),
    .in_id2_s_read(out_id_53__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_18__ap_start),
    .ap_done(krnl_globalSort_L1_L2_18__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_18__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_18__ap_ready),
    .in_dist0_s_dout(L1_out_dist_0__dout),
    .in_dist0_peek_dout(L1_out_dist_0__dout),
    .in_dist0_s_empty_n(L1_out_dist_0__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_0__empty_n),
    .in_dist0_s_read(L1_out_dist_0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_1__dout),
    .in_dist1_peek_dout(L1_out_dist_1__dout),
    .in_dist1_s_empty_n(L1_out_dist_1__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_1__empty_n),
    .in_dist1_s_read(L1_out_dist_1__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_2__dout),
    .in_dist2_peek_dout(L1_out_dist_2__dout),
    .in_dist2_s_empty_n(L1_out_dist_2__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_2__empty_n),
    .in_dist2_s_read(L1_out_dist_2__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_0__dout),
    .in_id0_peek_dout(L1_out_id_0__dout),
    .in_id0_s_empty_n(L1_out_id_0__empty_n),
    .in_id0_peek_empty_n(L1_out_id_0__empty_n),
    .in_id0_s_read(L1_out_id_0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_1__dout),
    .in_id1_peek_dout(L1_out_id_1__dout),
    .in_id1_s_empty_n(L1_out_id_1__empty_n),
    .in_id1_peek_empty_n(L1_out_id_1__empty_n),
    .in_id1_s_read(L1_out_id_1__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_2__dout),
    .in_id2_peek_dout(L1_out_id_2__dout),
    .in_id2_s_empty_n(L1_out_id_2__empty_n),
    .in_id2_peek_empty_n(L1_out_id_2__empty_n),
    .in_id2_s_read(L1_out_id_2__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist0__din),
    .out_dist_full_n(L2_out_dist0__full_n),
    .out_dist_write(L2_out_dist0__write),
    .out_id_din(L2_out_id0__din),
    .out_id_full_n(L2_out_id0__full_n),
    .out_id_write(L2_out_id0__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_19__ap_start),
    .ap_done(krnl_globalSort_L1_L2_19__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_19__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_19__ap_ready),
    .in_dist0_s_dout(L1_out_dist_3__dout),
    .in_dist0_peek_dout(L1_out_dist_3__dout),
    .in_dist0_s_empty_n(L1_out_dist_3__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_3__empty_n),
    .in_dist0_s_read(L1_out_dist_3__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_4__dout),
    .in_dist1_peek_dout(L1_out_dist_4__dout),
    .in_dist1_s_empty_n(L1_out_dist_4__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_4__empty_n),
    .in_dist1_s_read(L1_out_dist_4__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_5__dout),
    .in_dist2_peek_dout(L1_out_dist_5__dout),
    .in_dist2_s_empty_n(L1_out_dist_5__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_5__empty_n),
    .in_dist2_s_read(L1_out_dist_5__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_3__dout),
    .in_id0_peek_dout(L1_out_id_3__dout),
    .in_id0_s_empty_n(L1_out_id_3__empty_n),
    .in_id0_peek_empty_n(L1_out_id_3__empty_n),
    .in_id0_s_read(L1_out_id_3__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_4__dout),
    .in_id1_peek_dout(L1_out_id_4__dout),
    .in_id1_s_empty_n(L1_out_id_4__empty_n),
    .in_id1_peek_empty_n(L1_out_id_4__empty_n),
    .in_id1_s_read(L1_out_id_4__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_5__dout),
    .in_id2_peek_dout(L1_out_id_5__dout),
    .in_id2_s_empty_n(L1_out_id_5__empty_n),
    .in_id2_peek_empty_n(L1_out_id_5__empty_n),
    .in_id2_s_read(L1_out_id_5__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist1__din),
    .out_dist_full_n(L2_out_dist1__full_n),
    .out_dist_write(L2_out_dist1__write),
    .out_id_din(L2_out_id1__din),
    .out_id_full_n(L2_out_id1__full_n),
    .out_id_write(L2_out_id1__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_20__ap_start),
    .ap_done(krnl_globalSort_L1_L2_20__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_20__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_20__ap_ready),
    .in_dist0_s_dout(L1_out_dist_6__dout),
    .in_dist0_peek_dout(L1_out_dist_6__dout),
    .in_dist0_s_empty_n(L1_out_dist_6__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_6__empty_n),
    .in_dist0_s_read(L1_out_dist_6__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_7__dout),
    .in_dist1_peek_dout(L1_out_dist_7__dout),
    .in_dist1_s_empty_n(L1_out_dist_7__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_7__empty_n),
    .in_dist1_s_read(L1_out_dist_7__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_8__dout),
    .in_dist2_peek_dout(L1_out_dist_8__dout),
    .in_dist2_s_empty_n(L1_out_dist_8__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_8__empty_n),
    .in_dist2_s_read(L1_out_dist_8__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_6__dout),
    .in_id0_peek_dout(L1_out_id_6__dout),
    .in_id0_s_empty_n(L1_out_id_6__empty_n),
    .in_id0_peek_empty_n(L1_out_id_6__empty_n),
    .in_id0_s_read(L1_out_id_6__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_7__dout),
    .in_id1_peek_dout(L1_out_id_7__dout),
    .in_id1_s_empty_n(L1_out_id_7__empty_n),
    .in_id1_peek_empty_n(L1_out_id_7__empty_n),
    .in_id1_s_read(L1_out_id_7__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_8__dout),
    .in_id2_peek_dout(L1_out_id_8__dout),
    .in_id2_s_empty_n(L1_out_id_8__empty_n),
    .in_id2_peek_empty_n(L1_out_id_8__empty_n),
    .in_id2_s_read(L1_out_id_8__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist2__din),
    .out_dist_full_n(L2_out_dist2__full_n),
    .out_dist_write(L2_out_dist2__write),
    .out_id_din(L2_out_id2__din),
    .out_id_full_n(L2_out_id2__full_n),
    .out_id_write(L2_out_id2__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_21__ap_start),
    .ap_done(krnl_globalSort_L1_L2_21__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_21__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_21__ap_ready),
    .in_dist1_s_dout(L1_out_dist_10__dout),
    .in_dist1_peek_dout(L1_out_dist_10__dout),
    .in_dist1_s_empty_n(L1_out_dist_10__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_10__empty_n),
    .in_dist1_s_read(L1_out_dist_10__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_11__dout),
    .in_dist2_peek_dout(L1_out_dist_11__dout),
    .in_dist2_s_empty_n(L1_out_dist_11__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_11__empty_n),
    .in_dist2_s_read(L1_out_dist_11__read),
    .in_dist2_peek_read(),
    .in_dist0_s_dout(L1_out_dist_9__dout),
    .in_dist0_peek_dout(L1_out_dist_9__dout),
    .in_dist0_s_empty_n(L1_out_dist_9__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_9__empty_n),
    .in_dist0_s_read(L1_out_dist_9__read),
    .in_dist0_peek_read(),
    .in_id1_s_dout(L1_out_id_10__dout),
    .in_id1_peek_dout(L1_out_id_10__dout),
    .in_id1_s_empty_n(L1_out_id_10__empty_n),
    .in_id1_peek_empty_n(L1_out_id_10__empty_n),
    .in_id1_s_read(L1_out_id_10__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_11__dout),
    .in_id2_peek_dout(L1_out_id_11__dout),
    .in_id2_s_empty_n(L1_out_id_11__empty_n),
    .in_id2_peek_empty_n(L1_out_id_11__empty_n),
    .in_id2_s_read(L1_out_id_11__read),
    .in_id2_peek_read(),
    .in_id0_s_dout(L1_out_id_9__dout),
    .in_id0_peek_dout(L1_out_id_9__dout),
    .in_id0_s_empty_n(L1_out_id_9__empty_n),
    .in_id0_peek_empty_n(L1_out_id_9__empty_n),
    .in_id0_s_read(L1_out_id_9__read),
    .in_id0_peek_read(),
    .out_dist_din(L2_out_dist3__din),
    .out_dist_full_n(L2_out_dist3__full_n),
    .out_dist_write(L2_out_dist3__write),
    .out_id_din(L2_out_id3__din),
    .out_id_full_n(L2_out_id3__full_n),
    .out_id_write(L2_out_id3__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_22__ap_start),
    .ap_done(krnl_globalSort_L1_L2_22__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_22__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_22__ap_ready),
    .in_dist0_s_dout(L1_out_dist_12__dout),
    .in_dist0_peek_dout(L1_out_dist_12__dout),
    .in_dist0_s_empty_n(L1_out_dist_12__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_12__empty_n),
    .in_dist0_s_read(L1_out_dist_12__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_13__dout),
    .in_dist1_peek_dout(L1_out_dist_13__dout),
    .in_dist1_s_empty_n(L1_out_dist_13__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_13__empty_n),
    .in_dist1_s_read(L1_out_dist_13__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_14__dout),
    .in_dist2_peek_dout(L1_out_dist_14__dout),
    .in_dist2_s_empty_n(L1_out_dist_14__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_14__empty_n),
    .in_dist2_s_read(L1_out_dist_14__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_12__dout),
    .in_id0_peek_dout(L1_out_id_12__dout),
    .in_id0_s_empty_n(L1_out_id_12__empty_n),
    .in_id0_peek_empty_n(L1_out_id_12__empty_n),
    .in_id0_s_read(L1_out_id_12__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_13__dout),
    .in_id1_peek_dout(L1_out_id_13__dout),
    .in_id1_s_empty_n(L1_out_id_13__empty_n),
    .in_id1_peek_empty_n(L1_out_id_13__empty_n),
    .in_id1_s_read(L1_out_id_13__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_14__dout),
    .in_id2_peek_dout(L1_out_id_14__dout),
    .in_id2_s_empty_n(L1_out_id_14__empty_n),
    .in_id2_peek_empty_n(L1_out_id_14__empty_n),
    .in_id2_s_read(L1_out_id_14__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist4__din),
    .out_dist_full_n(L2_out_dist4__full_n),
    .out_dist_write(L2_out_dist4__write),
    .out_id_din(L2_out_id4__din),
    .out_id_full_n(L2_out_id4__full_n),
    .out_id_write(L2_out_id4__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_23__ap_start),
    .ap_done(krnl_globalSort_L1_L2_23__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_23__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_23__ap_ready),
    .in_dist0_s_dout(L1_out_dist_15__dout),
    .in_dist0_peek_dout(L1_out_dist_15__dout),
    .in_dist0_s_empty_n(L1_out_dist_15__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_15__empty_n),
    .in_dist0_s_read(L1_out_dist_15__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_16__dout),
    .in_dist1_peek_dout(L1_out_dist_16__dout),
    .in_dist1_s_empty_n(L1_out_dist_16__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_16__empty_n),
    .in_dist1_s_read(L1_out_dist_16__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_17__dout),
    .in_dist2_peek_dout(L1_out_dist_17__dout),
    .in_dist2_s_empty_n(L1_out_dist_17__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_17__empty_n),
    .in_dist2_s_read(L1_out_dist_17__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_15__dout),
    .in_id0_peek_dout(L1_out_id_15__dout),
    .in_id0_s_empty_n(L1_out_id_15__empty_n),
    .in_id0_peek_empty_n(L1_out_id_15__empty_n),
    .in_id0_s_read(L1_out_id_15__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_16__dout),
    .in_id1_peek_dout(L1_out_id_16__dout),
    .in_id1_s_empty_n(L1_out_id_16__empty_n),
    .in_id1_peek_empty_n(L1_out_id_16__empty_n),
    .in_id1_s_read(L1_out_id_16__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_17__dout),
    .in_id2_peek_dout(L1_out_id_17__dout),
    .in_id2_s_empty_n(L1_out_id_17__empty_n),
    .in_id2_peek_empty_n(L1_out_id_17__empty_n),
    .in_id2_s_read(L1_out_id_17__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist5__din),
    .out_dist_full_n(L2_out_dist5__full_n),
    .out_dist_write(L2_out_dist5__write),
    .out_id_din(L2_out_id5__din),
    .out_id_full_n(L2_out_id5__full_n),
    .out_id_write(L2_out_id5__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_24__ap_start),
    .ap_done(krnl_globalSort_L1_L2_24__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_24__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_24__ap_ready),
    .in_dist0_s_dout(L2_out_dist0__dout),
    .in_dist0_peek_dout(L2_out_dist0__dout),
    .in_dist0_s_empty_n(L2_out_dist0__empty_n),
    .in_dist0_peek_empty_n(L2_out_dist0__empty_n),
    .in_dist0_s_read(L2_out_dist0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L2_out_dist1__dout),
    .in_dist1_peek_dout(L2_out_dist1__dout),
    .in_dist1_s_empty_n(L2_out_dist1__empty_n),
    .in_dist1_peek_empty_n(L2_out_dist1__empty_n),
    .in_dist1_s_read(L2_out_dist1__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L2_out_dist2__dout),
    .in_dist2_peek_dout(L2_out_dist2__dout),
    .in_dist2_s_empty_n(L2_out_dist2__empty_n),
    .in_dist2_peek_empty_n(L2_out_dist2__empty_n),
    .in_dist2_s_read(L2_out_dist2__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L2_out_id0__dout),
    .in_id0_peek_dout(L2_out_id0__dout),
    .in_id0_s_empty_n(L2_out_id0__empty_n),
    .in_id0_peek_empty_n(L2_out_id0__empty_n),
    .in_id0_s_read(L2_out_id0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L2_out_id1__dout),
    .in_id1_peek_dout(L2_out_id1__dout),
    .in_id1_s_empty_n(L2_out_id1__empty_n),
    .in_id1_peek_empty_n(L2_out_id1__empty_n),
    .in_id1_s_read(L2_out_id1__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L2_out_id2__dout),
    .in_id2_peek_dout(L2_out_id2__dout),
    .in_id2_s_empty_n(L2_out_id2__empty_n),
    .in_id2_peek_empty_n(L2_out_id2__empty_n),
    .in_id2_s_read(L2_out_id2__read),
    .in_id2_peek_read(),
    .out_dist_din(L3_out_dist0__din),
    .out_dist_full_n(L3_out_dist0__full_n),
    .out_dist_write(L3_out_dist0__write),
    .out_id_din(L3_out_id0__din),
    .out_id_full_n(L3_out_id0__full_n),
    .out_id_write(L3_out_id0__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_25__ap_start),
    .ap_done(krnl_globalSort_L1_L2_25__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_25__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_25__ap_ready),
    .in_dist0_s_dout(L2_out_dist3__dout),
    .in_dist0_peek_dout(L2_out_dist3__dout),
    .in_dist0_s_empty_n(L2_out_dist3__empty_n),
    .in_dist0_peek_empty_n(L2_out_dist3__empty_n),
    .in_dist0_s_read(L2_out_dist3__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L2_out_dist4__dout),
    .in_dist1_peek_dout(L2_out_dist4__dout),
    .in_dist1_s_empty_n(L2_out_dist4__empty_n),
    .in_dist1_peek_empty_n(L2_out_dist4__empty_n),
    .in_dist1_s_read(L2_out_dist4__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L2_out_dist5__dout),
    .in_dist2_peek_dout(L2_out_dist5__dout),
    .in_dist2_s_empty_n(L2_out_dist5__empty_n),
    .in_dist2_peek_empty_n(L2_out_dist5__empty_n),
    .in_dist2_s_read(L2_out_dist5__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L2_out_id3__dout),
    .in_id0_peek_dout(L2_out_id3__dout),
    .in_id0_s_empty_n(L2_out_id3__empty_n),
    .in_id0_peek_empty_n(L2_out_id3__empty_n),
    .in_id0_s_read(L2_out_id3__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L2_out_id4__dout),
    .in_id1_peek_dout(L2_out_id4__dout),
    .in_id1_s_empty_n(L2_out_id4__empty_n),
    .in_id1_peek_empty_n(L2_out_id4__empty_n),
    .in_id1_s_read(L2_out_id4__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L2_out_id5__dout),
    .in_id2_peek_dout(L2_out_id5__dout),
    .in_id2_s_empty_n(L2_out_id5__empty_n),
    .in_id2_peek_empty_n(L2_out_id5__empty_n),
    .in_id2_s_read(L2_out_id5__read),
    .in_id2_peek_read(),
    .out_dist_din(L3_out_dist1__din),
    .out_dist_full_n(L3_out_dist1__full_n),
    .out_dist_write(L3_out_dist1__write),
    .out_id_din(L3_out_id1__din),
    .out_id_full_n(L3_out_id1__full_n),
    .out_id_write(L3_out_id1__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L3
  krnl_globalSort_L3_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L3_0__ap_start),
    .ap_done(krnl_globalSort_L3_0__ap_done),
    .ap_idle(krnl_globalSort_L3_0__ap_idle),
    .ap_ready(krnl_globalSort_L3_0__ap_ready),
    .in_dist0_s_dout(L3_out_dist0__dout),
    .in_dist0_peek_dout(L3_out_dist0__dout),
    .in_dist0_s_empty_n(L3_out_dist0__empty_n),
    .in_dist0_peek_empty_n(L3_out_dist0__empty_n),
    .in_dist0_s_read(L3_out_dist0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L3_out_dist1__dout),
    .in_dist1_peek_dout(L3_out_dist1__dout),
    .in_dist1_s_empty_n(L3_out_dist1__empty_n),
    .in_dist1_peek_empty_n(L3_out_dist1__empty_n),
    .in_dist1_s_read(L3_out_dist1__read),
    .in_dist1_peek_read(),
    .in_id0_s_dout(L3_out_id0__dout),
    .in_id0_peek_dout(L3_out_id0__dout),
    .in_id0_s_empty_n(L3_out_id0__empty_n),
    .in_id0_peek_empty_n(L3_out_id0__empty_n),
    .in_id0_s_read(L3_out_id0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L3_out_id1__dout),
    .in_id1_peek_dout(L3_out_id1__dout),
    .in_id1_s_empty_n(L3_out_id1__empty_n),
    .in_id1_peek_empty_n(L3_out_id1__empty_n),
    .in_id1_s_read(L3_out_id1__read),
    .in_id1_peek_read(),
    .output_knnDist_read_addr_s_din(L4_out_dist_read_addr__din),
    .output_knnDist_read_addr_s_full_n(L4_out_dist_read_addr__full_n),
    .output_knnDist_read_addr_s_write(L4_out_dist_read_addr__write),
    .output_knnDist_read_addr_offset(krnl_globalSort_L3_0___L4_out_dist__q0),
    .output_knnDist_read_data_s_dout({1'b0, L4_out_dist_read_data__dout}),
    .output_knnDist_read_data_peek_dout({1'b0, L4_out_dist_read_data__dout}),
    .output_knnDist_read_data_s_empty_n(L4_out_dist_read_data__empty_n),
    .output_knnDist_read_data_peek_empty_n(L4_out_dist_read_data__empty_n),
    .output_knnDist_read_data_s_read(L4_out_dist_read_data__read),
    .output_knnDist_read_data_peek_read(),
    .output_knnDist_write_addr_s_din(L4_out_dist_write_addr__din),
    .output_knnDist_write_addr_s_full_n(L4_out_dist_write_addr__full_n),
    .output_knnDist_write_addr_s_write(L4_out_dist_write_addr__write),
    .output_knnDist_write_addr_offset(krnl_globalSort_L3_0___L4_out_dist__q0),
    .output_knnDist_write_data_din(L4_out_dist_write_data__din),
    .output_knnDist_write_data_full_n(L4_out_dist_write_data__full_n),
    .output_knnDist_write_data_write(L4_out_dist_write_data__write),
    .output_knnDist_write_resp_s_dout({1'b0, L4_out_dist_write_resp__dout}),
    .output_knnDist_write_resp_peek_dout({1'b0, L4_out_dist_write_resp__dout}),
    .output_knnDist_write_resp_s_empty_n(L4_out_dist_write_resp__empty_n),
    .output_knnDist_write_resp_peek_empty_n(L4_out_dist_write_resp__empty_n),
    .output_knnDist_write_resp_s_read(L4_out_dist_write_resp__read),
    .output_knnDist_write_resp_peek_read(),
    .output_knnId_read_addr_s_din(L4_out_id_read_addr__din),
    .output_knnId_read_addr_s_full_n(L4_out_id_read_addr__full_n),
    .output_knnId_read_addr_s_write(L4_out_id_read_addr__write),
    .output_knnId_read_addr_offset(krnl_globalSort_L3_0___L4_out_id__q0),
    .output_knnId_read_data_s_dout({1'b0, L4_out_id_read_data__dout}),
    .output_knnId_read_data_peek_dout({1'b0, L4_out_id_read_data__dout}),
    .output_knnId_read_data_s_empty_n(L4_out_id_read_data__empty_n),
    .output_knnId_read_data_peek_empty_n(L4_out_id_read_data__empty_n),
    .output_knnId_read_data_s_read(L4_out_id_read_data__read),
    .output_knnId_read_data_peek_read(),
    .output_knnId_write_addr_s_din(L4_out_id_write_addr__din),
    .output_knnId_write_addr_s_full_n(L4_out_id_write_addr__full_n),
    .output_knnId_write_addr_s_write(L4_out_id_write_addr__write),
    .output_knnId_write_addr_offset(krnl_globalSort_L3_0___L4_out_id__q0),
    .output_knnId_write_data_din(L4_out_id_write_data__din),
    .output_knnId_write_data_full_n(L4_out_id_write_data__full_n),
    .output_knnId_write_data_write(L4_out_id_write_data__write),
    .output_knnId_write_resp_s_dout({1'b0, L4_out_id_write_resp__dout}),
    .output_knnId_write_resp_peek_dout({1'b0, L4_out_id_write_resp__dout}),
    .output_knnId_write_resp_s_empty_n(L4_out_id_write_resp__empty_n),
    .output_knnId_write_resp_peek_empty_n(L4_out_id_write_resp__empty_n),
    .output_knnId_write_resp_s_read(L4_out_id_write_resp__read),
    .output_knnId_write_resp_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_0
  krnl_partialKnn_wrapper_0_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_0_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_0_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_0_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_0_0__ap_ready),
    .start_id_0(64'd0),
    .searchSpace_0_read_addr_s_din(in_0_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_0_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_0_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_0_0___in_0__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_0_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_0_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_0_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_0_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_0_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_0_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_0_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_0_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_0_0___in_0__q0),
    .searchSpace_0_write_data_din(in_0_write_data__din),
    .searchSpace_0_write_data_full_n(in_0_write_data__full_n),
    .searchSpace_0_write_data_write(in_0_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_0_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_0_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_0_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_0_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_0_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_0__din),
    .out_dist_full_n(out_dist_0__full_n),
    .out_dist_write(out_dist_0__write),
    .out_id_din(out_id_0__din),
    .out_id_full_n(out_id_0__full_n),
    .out_id_write(out_id_0__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_1
  krnl_partialKnn_wrapper_1_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_1_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_1_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_1_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_1_0__ap_ready),
    .start_id_0(64'd8192),
    .searchSpace_0_read_addr_s_din(in_1_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_1_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_1_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_1_0___in_1__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_1_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_1_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_1_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_1_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_1_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_1_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_1_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_1_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_1_0___in_1__q0),
    .searchSpace_0_write_data_din(in_1_write_data__din),
    .searchSpace_0_write_data_full_n(in_1_write_data__full_n),
    .searchSpace_0_write_data_write(in_1_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_1_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_1_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_1_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_1_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_1_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_1__din),
    .out_dist_full_n(out_dist_1__full_n),
    .out_dist_write(out_dist_1__write),
    .out_id_din(out_id_1__din),
    .out_id_full_n(out_id_1__full_n),
    .out_id_write(out_id_1__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_10
  krnl_partialKnn_wrapper_10_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_10_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_10_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_10_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_10_0__ap_ready),
    .start_id_0(64'd81920),
    .searchSpace_0_read_addr_s_din(in_10_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_10_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_10_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_10_0___in_10__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_10_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_10_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_10_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_10_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_10_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_10_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_10_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_10_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_10_0___in_10__q0),
    .searchSpace_0_write_data_din(in_10_write_data__din),
    .searchSpace_0_write_data_full_n(in_10_write_data__full_n),
    .searchSpace_0_write_data_write(in_10_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_10_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_10_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_10_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_10_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_10_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_10__din),
    .out_dist_full_n(out_dist_10__full_n),
    .out_dist_write(out_dist_10__write),
    .out_id_din(out_id_10__din),
    .out_id_full_n(out_id_10__full_n),
    .out_id_write(out_id_10__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_11
  krnl_partialKnn_wrapper_11_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_11_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_11_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_11_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_11_0__ap_ready),
    .start_id_0(64'd90112),
    .searchSpace_0_read_addr_s_din(in_11_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_11_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_11_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_11_0___in_11__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_11_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_11_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_11_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_11_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_11_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_11_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_11_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_11_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_11_0___in_11__q0),
    .searchSpace_0_write_data_din(in_11_write_data__din),
    .searchSpace_0_write_data_full_n(in_11_write_data__full_n),
    .searchSpace_0_write_data_write(in_11_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_11_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_11_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_11_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_11_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_11_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_11__din),
    .out_dist_full_n(out_dist_11__full_n),
    .out_dist_write(out_dist_11__write),
    .out_id_din(out_id_11__din),
    .out_id_full_n(out_id_11__full_n),
    .out_id_write(out_id_11__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_12
  krnl_partialKnn_wrapper_12_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_12_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_12_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_12_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_12_0__ap_ready),
    .start_id_0(64'd98304),
    .searchSpace_0_read_addr_s_din(in_12_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_12_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_12_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_12_0___in_12__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_12_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_12_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_12_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_12_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_12_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_12_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_12_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_12_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_12_0___in_12__q0),
    .searchSpace_0_write_data_din(in_12_write_data__din),
    .searchSpace_0_write_data_full_n(in_12_write_data__full_n),
    .searchSpace_0_write_data_write(in_12_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_12_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_12_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_12_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_12_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_12_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_12__din),
    .out_dist_full_n(out_dist_12__full_n),
    .out_dist_write(out_dist_12__write),
    .out_id_din(out_id_12__din),
    .out_id_full_n(out_id_12__full_n),
    .out_id_write(out_id_12__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_13
  krnl_partialKnn_wrapper_13_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_13_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_13_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_13_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_13_0__ap_ready),
    .start_id_0(64'd106496),
    .searchSpace_0_read_addr_s_din(in_13_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_13_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_13_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_13_0___in_13__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_13_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_13_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_13_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_13_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_13_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_13_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_13_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_13_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_13_0___in_13__q0),
    .searchSpace_0_write_data_din(in_13_write_data__din),
    .searchSpace_0_write_data_full_n(in_13_write_data__full_n),
    .searchSpace_0_write_data_write(in_13_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_13_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_13_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_13_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_13_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_13_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_13__din),
    .out_dist_full_n(out_dist_13__full_n),
    .out_dist_write(out_dist_13__write),
    .out_id_din(out_id_13__din),
    .out_id_full_n(out_id_13__full_n),
    .out_id_write(out_id_13__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_14
  krnl_partialKnn_wrapper_14_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_14_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_14_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_14_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_14_0__ap_ready),
    .start_id_0(64'd114688),
    .searchSpace_0_read_addr_s_din(in_14_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_14_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_14_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_14_0___in_14__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_14_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_14_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_14_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_14_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_14_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_14_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_14_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_14_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_14_0___in_14__q0),
    .searchSpace_0_write_data_din(in_14_write_data__din),
    .searchSpace_0_write_data_full_n(in_14_write_data__full_n),
    .searchSpace_0_write_data_write(in_14_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_14_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_14_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_14_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_14_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_14_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_14__din),
    .out_dist_full_n(out_dist_14__full_n),
    .out_dist_write(out_dist_14__write),
    .out_id_din(out_id_14__din),
    .out_id_full_n(out_id_14__full_n),
    .out_id_write(out_id_14__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_15
  krnl_partialKnn_wrapper_15_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_15_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_15_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_15_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_15_0__ap_ready),
    .start_id_0(64'd122880),
    .searchSpace_0_read_addr_s_din(in_15_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_15_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_15_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_15_0___in_15__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_15_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_15_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_15_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_15_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_15_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_15_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_15_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_15_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_15_0___in_15__q0),
    .searchSpace_0_write_data_din(in_15_write_data__din),
    .searchSpace_0_write_data_full_n(in_15_write_data__full_n),
    .searchSpace_0_write_data_write(in_15_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_15_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_15_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_15_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_15_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_15_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_15__din),
    .out_dist_full_n(out_dist_15__full_n),
    .out_dist_write(out_dist_15__write),
    .out_id_din(out_id_15__din),
    .out_id_full_n(out_id_15__full_n),
    .out_id_write(out_id_15__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_16
  krnl_partialKnn_wrapper_16_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_16_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_16_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_16_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_16_0__ap_ready),
    .start_id_0(64'd131072),
    .searchSpace_0_read_addr_s_din(in_16_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_16_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_16_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_16_0___in_16__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_16_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_16_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_16_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_16_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_16_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_16_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_16_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_16_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_16_0___in_16__q0),
    .searchSpace_0_write_data_din(in_16_write_data__din),
    .searchSpace_0_write_data_full_n(in_16_write_data__full_n),
    .searchSpace_0_write_data_write(in_16_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_16_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_16_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_16_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_16_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_16_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_16__din),
    .out_dist_full_n(out_dist_16__full_n),
    .out_dist_write(out_dist_16__write),
    .out_id_din(out_id_16__din),
    .out_id_full_n(out_id_16__full_n),
    .out_id_write(out_id_16__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_17
  krnl_partialKnn_wrapper_17_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_17_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_17_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_17_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_17_0__ap_ready),
    .start_id_0(64'd139264),
    .searchSpace_0_read_addr_s_din(in_17_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_17_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_17_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_17_0___in_17__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_17_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_17_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_17_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_17_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_17_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_17_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_17_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_17_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_17_0___in_17__q0),
    .searchSpace_0_write_data_din(in_17_write_data__din),
    .searchSpace_0_write_data_full_n(in_17_write_data__full_n),
    .searchSpace_0_write_data_write(in_17_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_17_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_17_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_17_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_17_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_17_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_17__din),
    .out_dist_full_n(out_dist_17__full_n),
    .out_dist_write(out_dist_17__write),
    .out_id_din(out_id_17__din),
    .out_id_full_n(out_id_17__full_n),
    .out_id_write(out_id_17__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_18
  krnl_partialKnn_wrapper_18_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_18_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_18_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_18_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_18_0__ap_ready),
    .start_id_0(64'd147456),
    .searchSpace_0_read_addr_s_din(in_18_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_18_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_18_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_18_0___in_18__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_18_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_18_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_18_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_18_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_18_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_18_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_18_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_18_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_18_0___in_18__q0),
    .searchSpace_0_write_data_din(in_18_write_data__din),
    .searchSpace_0_write_data_full_n(in_18_write_data__full_n),
    .searchSpace_0_write_data_write(in_18_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_18_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_18_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_18_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_18_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_18_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_18__din),
    .out_dist_full_n(out_dist_18__full_n),
    .out_dist_write(out_dist_18__write),
    .out_id_din(out_id_18__din),
    .out_id_full_n(out_id_18__full_n),
    .out_id_write(out_id_18__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_19
  krnl_partialKnn_wrapper_19_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_19_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_19_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_19_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_19_0__ap_ready),
    .start_id_0(64'd155648),
    .searchSpace_0_read_addr_s_din(in_19_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_19_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_19_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_19_0___in_19__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_19_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_19_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_19_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_19_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_19_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_19_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_19_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_19_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_19_0___in_19__q0),
    .searchSpace_0_write_data_din(in_19_write_data__din),
    .searchSpace_0_write_data_full_n(in_19_write_data__full_n),
    .searchSpace_0_write_data_write(in_19_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_19_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_19_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_19_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_19_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_19_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_19__din),
    .out_dist_full_n(out_dist_19__full_n),
    .out_dist_write(out_dist_19__write),
    .out_id_din(out_id_19__din),
    .out_id_full_n(out_id_19__full_n),
    .out_id_write(out_id_19__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_2
  krnl_partialKnn_wrapper_2_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_2_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_2_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_2_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_2_0__ap_ready),
    .start_id_0(64'd16384),
    .searchSpace_0_read_addr_s_din(in_2_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_2_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_2_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_2_0___in_2__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_2_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_2_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_2_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_2_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_2_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_2_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_2_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_2_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_2_0___in_2__q0),
    .searchSpace_0_write_data_din(in_2_write_data__din),
    .searchSpace_0_write_data_full_n(in_2_write_data__full_n),
    .searchSpace_0_write_data_write(in_2_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_2_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_2_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_2_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_2_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_2_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_2__din),
    .out_dist_full_n(out_dist_2__full_n),
    .out_dist_write(out_dist_2__write),
    .out_id_din(out_id_2__din),
    .out_id_full_n(out_id_2__full_n),
    .out_id_write(out_id_2__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_20
  krnl_partialKnn_wrapper_20_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_20_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_20_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_20_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_20_0__ap_ready),
    .start_id_0(64'd163840),
    .searchSpace_0_read_addr_s_din(in_20_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_20_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_20_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_20_0___in_20__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_20_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_20_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_20_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_20_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_20_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_20_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_20_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_20_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_20_0___in_20__q0),
    .searchSpace_0_write_data_din(in_20_write_data__din),
    .searchSpace_0_write_data_full_n(in_20_write_data__full_n),
    .searchSpace_0_write_data_write(in_20_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_20_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_20_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_20_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_20_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_20_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_20__din),
    .out_dist_full_n(out_dist_20__full_n),
    .out_dist_write(out_dist_20__write),
    .out_id_din(out_id_20__din),
    .out_id_full_n(out_id_20__full_n),
    .out_id_write(out_id_20__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_21
  krnl_partialKnn_wrapper_21_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_21_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_21_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_21_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_21_0__ap_ready),
    .start_id_0(64'd172032),
    .searchSpace_0_read_addr_s_din(in_21_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_21_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_21_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_21_0___in_21__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_21_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_21_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_21_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_21_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_21_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_21_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_21_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_21_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_21_0___in_21__q0),
    .searchSpace_0_write_data_din(in_21_write_data__din),
    .searchSpace_0_write_data_full_n(in_21_write_data__full_n),
    .searchSpace_0_write_data_write(in_21_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_21_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_21_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_21_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_21_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_21_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_21__din),
    .out_dist_full_n(out_dist_21__full_n),
    .out_dist_write(out_dist_21__write),
    .out_id_din(out_id_21__din),
    .out_id_full_n(out_id_21__full_n),
    .out_id_write(out_id_21__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_22
  krnl_partialKnn_wrapper_22_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_22_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_22_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_22_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_22_0__ap_ready),
    .start_id_0(64'd180224),
    .searchSpace_0_read_addr_s_din(in_22_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_22_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_22_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_22_0___in_22__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_22_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_22_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_22_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_22_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_22_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_22_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_22_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_22_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_22_0___in_22__q0),
    .searchSpace_0_write_data_din(in_22_write_data__din),
    .searchSpace_0_write_data_full_n(in_22_write_data__full_n),
    .searchSpace_0_write_data_write(in_22_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_22_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_22_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_22_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_22_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_22_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_22__din),
    .out_dist_full_n(out_dist_22__full_n),
    .out_dist_write(out_dist_22__write),
    .out_id_din(out_id_22__din),
    .out_id_full_n(out_id_22__full_n),
    .out_id_write(out_id_22__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_23
  krnl_partialKnn_wrapper_23_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_23_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_23_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_23_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_23_0__ap_ready),
    .start_id_0(64'd188416),
    .searchSpace_0_read_addr_s_din(in_23_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_23_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_23_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_23_0___in_23__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_23_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_23_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_23_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_23_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_23_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_23_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_23_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_23_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_23_0___in_23__q0),
    .searchSpace_0_write_data_din(in_23_write_data__din),
    .searchSpace_0_write_data_full_n(in_23_write_data__full_n),
    .searchSpace_0_write_data_write(in_23_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_23_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_23_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_23_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_23_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_23_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_23__din),
    .out_dist_full_n(out_dist_23__full_n),
    .out_dist_write(out_dist_23__write),
    .out_id_din(out_id_23__din),
    .out_id_full_n(out_id_23__full_n),
    .out_id_write(out_id_23__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_24
  krnl_partialKnn_wrapper_24_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_24_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_24_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_24_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_24_0__ap_ready),
    .start_id_0(64'd196608),
    .searchSpace_0_read_addr_s_din(in_24_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_24_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_24_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_24_0___in_24__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_24_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_24_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_24_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_24_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_24_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_24_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_24_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_24_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_24_0___in_24__q0),
    .searchSpace_0_write_data_din(in_24_write_data__din),
    .searchSpace_0_write_data_full_n(in_24_write_data__full_n),
    .searchSpace_0_write_data_write(in_24_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_24_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_24_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_24_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_24_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_24_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_24__din),
    .out_dist_full_n(out_dist_24__full_n),
    .out_dist_write(out_dist_24__write),
    .out_id_din(out_id_24__din),
    .out_id_full_n(out_id_24__full_n),
    .out_id_write(out_id_24__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_25
  krnl_partialKnn_wrapper_25_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_25_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_25_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_25_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_25_0__ap_ready),
    .start_id_0(64'd204800),
    .searchSpace_0_read_addr_s_din(in_25_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_25_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_25_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_25_0___in_25__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_25_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_25_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_25_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_25_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_25_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_25_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_25_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_25_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_25_0___in_25__q0),
    .searchSpace_0_write_data_din(in_25_write_data__din),
    .searchSpace_0_write_data_full_n(in_25_write_data__full_n),
    .searchSpace_0_write_data_write(in_25_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_25_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_25_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_25_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_25_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_25_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_25__din),
    .out_dist_full_n(out_dist_25__full_n),
    .out_dist_write(out_dist_25__write),
    .out_id_din(out_id_25__din),
    .out_id_full_n(out_id_25__full_n),
    .out_id_write(out_id_25__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_26
  krnl_partialKnn_wrapper_26_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_26_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_26_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_26_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_26_0__ap_ready),
    .start_id_0(64'd212992),
    .searchSpace_0_read_addr_s_din(in_26_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_26_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_26_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_26_0___in_26__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_26_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_26_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_26_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_26_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_26_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_26_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_26_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_26_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_26_0___in_26__q0),
    .searchSpace_0_write_data_din(in_26_write_data__din),
    .searchSpace_0_write_data_full_n(in_26_write_data__full_n),
    .searchSpace_0_write_data_write(in_26_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_26_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_26_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_26_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_26_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_26_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_26__din),
    .out_dist_full_n(out_dist_26__full_n),
    .out_dist_write(out_dist_26__write),
    .out_id_din(out_id_26__din),
    .out_id_full_n(out_id_26__full_n),
    .out_id_write(out_id_26__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_27
  krnl_partialKnn_wrapper_27_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_27_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_27_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_27_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_27_0__ap_ready),
    .start_id_0(64'd221184),
    .searchSpace_0_read_addr_s_din(in_27_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_27_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_27_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_27_0___in_27__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_27_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_27_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_27_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_27_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_27_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_27_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_27_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_27_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_27_0___in_27__q0),
    .searchSpace_0_write_data_din(in_27_write_data__din),
    .searchSpace_0_write_data_full_n(in_27_write_data__full_n),
    .searchSpace_0_write_data_write(in_27_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_27_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_27_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_27_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_27_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_27_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_27__din),
    .out_dist_full_n(out_dist_27__full_n),
    .out_dist_write(out_dist_27__write),
    .out_id_din(out_id_27__din),
    .out_id_full_n(out_id_27__full_n),
    .out_id_write(out_id_27__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_28
  krnl_partialKnn_wrapper_28_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_28_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_28_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_28_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_28_0__ap_ready),
    .start_id_0(64'd229376),
    .searchSpace_0_read_addr_s_din(in_28_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_28_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_28_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_28_0___in_28__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_28_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_28_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_28_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_28_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_28_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_28_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_28_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_28_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_28_0___in_28__q0),
    .searchSpace_0_write_data_din(in_28_write_data__din),
    .searchSpace_0_write_data_full_n(in_28_write_data__full_n),
    .searchSpace_0_write_data_write(in_28_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_28_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_28_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_28_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_28_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_28_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_28__din),
    .out_dist_full_n(out_dist_28__full_n),
    .out_dist_write(out_dist_28__write),
    .out_id_din(out_id_28__din),
    .out_id_full_n(out_id_28__full_n),
    .out_id_write(out_id_28__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_29
  krnl_partialKnn_wrapper_29_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_29_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_29_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_29_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_29_0__ap_ready),
    .start_id_0(64'd237568),
    .searchSpace_0_read_addr_s_din(in_29_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_29_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_29_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_29_0___in_29__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_29_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_29_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_29_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_29_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_29_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_29_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_29_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_29_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_29_0___in_29__q0),
    .searchSpace_0_write_data_din(in_29_write_data__din),
    .searchSpace_0_write_data_full_n(in_29_write_data__full_n),
    .searchSpace_0_write_data_write(in_29_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_29_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_29_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_29_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_29_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_29_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_29__din),
    .out_dist_full_n(out_dist_29__full_n),
    .out_dist_write(out_dist_29__write),
    .out_id_din(out_id_29__din),
    .out_id_full_n(out_id_29__full_n),
    .out_id_write(out_id_29__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_3
  krnl_partialKnn_wrapper_3_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_3_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_3_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_3_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_3_0__ap_ready),
    .start_id_0(64'd24576),
    .searchSpace_0_read_addr_s_din(in_3_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_3_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_3_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_3_0___in_3__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_3_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_3_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_3_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_3_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_3_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_3_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_3_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_3_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_3_0___in_3__q0),
    .searchSpace_0_write_data_din(in_3_write_data__din),
    .searchSpace_0_write_data_full_n(in_3_write_data__full_n),
    .searchSpace_0_write_data_write(in_3_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_3_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_3_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_3_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_3_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_3_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_3__din),
    .out_dist_full_n(out_dist_3__full_n),
    .out_dist_write(out_dist_3__write),
    .out_id_din(out_id_3__din),
    .out_id_full_n(out_id_3__full_n),
    .out_id_write(out_id_3__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_30
  krnl_partialKnn_wrapper_30_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_30_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_30_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_30_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_30_0__ap_ready),
    .start_id_0(64'd245760),
    .searchSpace_0_read_addr_s_din(in_30_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_30_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_30_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_30_0___in_30__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_30_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_30_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_30_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_30_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_30_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_30_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_30_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_30_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_30_0___in_30__q0),
    .searchSpace_0_write_data_din(in_30_write_data__din),
    .searchSpace_0_write_data_full_n(in_30_write_data__full_n),
    .searchSpace_0_write_data_write(in_30_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_30_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_30_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_30_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_30_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_30_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_30__din),
    .out_dist_full_n(out_dist_30__full_n),
    .out_dist_write(out_dist_30__write),
    .out_id_din(out_id_30__din),
    .out_id_full_n(out_id_30__full_n),
    .out_id_write(out_id_30__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_31
  krnl_partialKnn_wrapper_31_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_31_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_31_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_31_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_31_0__ap_ready),
    .start_id_0(64'd253952),
    .searchSpace_0_read_addr_s_din(in_31_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_31_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_31_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_31_0___in_31__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_31_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_31_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_31_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_31_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_31_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_31_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_31_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_31_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_31_0___in_31__q0),
    .searchSpace_0_write_data_din(in_31_write_data__din),
    .searchSpace_0_write_data_full_n(in_31_write_data__full_n),
    .searchSpace_0_write_data_write(in_31_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_31_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_31_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_31_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_31_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_31_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_31__din),
    .out_dist_full_n(out_dist_31__full_n),
    .out_dist_write(out_dist_31__write),
    .out_id_din(out_id_31__din),
    .out_id_full_n(out_id_31__full_n),
    .out_id_write(out_id_31__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_32
  krnl_partialKnn_wrapper_32_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_32_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_32_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_32_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_32_0__ap_ready),
    .start_id_0(64'd262144),
    .searchSpace_0_read_addr_s_din(in_32_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_32_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_32_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_32_0___in_32__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_32_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_32_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_32_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_32_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_32_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_32_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_32_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_32_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_32_0___in_32__q0),
    .searchSpace_0_write_data_din(in_32_write_data__din),
    .searchSpace_0_write_data_full_n(in_32_write_data__full_n),
    .searchSpace_0_write_data_write(in_32_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_32_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_32_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_32_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_32_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_32_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_32__din),
    .out_dist_full_n(out_dist_32__full_n),
    .out_dist_write(out_dist_32__write),
    .out_id_din(out_id_32__din),
    .out_id_full_n(out_id_32__full_n),
    .out_id_write(out_id_32__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_33
  krnl_partialKnn_wrapper_33_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_33_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_33_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_33_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_33_0__ap_ready),
    .start_id_0(64'd270336),
    .searchSpace_0_read_addr_s_din(in_33_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_33_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_33_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_33_0___in_33__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_33_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_33_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_33_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_33_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_33_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_33_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_33_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_33_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_33_0___in_33__q0),
    .searchSpace_0_write_data_din(in_33_write_data__din),
    .searchSpace_0_write_data_full_n(in_33_write_data__full_n),
    .searchSpace_0_write_data_write(in_33_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_33_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_33_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_33_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_33_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_33_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_33__din),
    .out_dist_full_n(out_dist_33__full_n),
    .out_dist_write(out_dist_33__write),
    .out_id_din(out_id_33__din),
    .out_id_full_n(out_id_33__full_n),
    .out_id_write(out_id_33__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_34
  krnl_partialKnn_wrapper_34_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_34_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_34_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_34_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_34_0__ap_ready),
    .start_id_0(64'd278528),
    .searchSpace_0_read_addr_s_din(in_34_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_34_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_34_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_34_0___in_34__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_34_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_34_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_34_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_34_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_34_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_34_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_34_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_34_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_34_0___in_34__q0),
    .searchSpace_0_write_data_din(in_34_write_data__din),
    .searchSpace_0_write_data_full_n(in_34_write_data__full_n),
    .searchSpace_0_write_data_write(in_34_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_34_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_34_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_34_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_34_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_34_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_34__din),
    .out_dist_full_n(out_dist_34__full_n),
    .out_dist_write(out_dist_34__write),
    .out_id_din(out_id_34__din),
    .out_id_full_n(out_id_34__full_n),
    .out_id_write(out_id_34__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_35
  krnl_partialKnn_wrapper_35_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_35_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_35_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_35_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_35_0__ap_ready),
    .start_id_0(64'd286720),
    .searchSpace_0_read_addr_s_din(in_35_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_35_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_35_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_35_0___in_35__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_35_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_35_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_35_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_35_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_35_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_35_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_35_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_35_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_35_0___in_35__q0),
    .searchSpace_0_write_data_din(in_35_write_data__din),
    .searchSpace_0_write_data_full_n(in_35_write_data__full_n),
    .searchSpace_0_write_data_write(in_35_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_35_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_35_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_35_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_35_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_35_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_35__din),
    .out_dist_full_n(out_dist_35__full_n),
    .out_dist_write(out_dist_35__write),
    .out_id_din(out_id_35__din),
    .out_id_full_n(out_id_35__full_n),
    .out_id_write(out_id_35__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_36
  krnl_partialKnn_wrapper_36_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_36_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_36_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_36_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_36_0__ap_ready),
    .start_id_0(64'd294912),
    .searchSpace_0_read_addr_s_din(in_36_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_36_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_36_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_36_0___in_36__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_36_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_36_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_36_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_36_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_36_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_36_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_36_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_36_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_36_0___in_36__q0),
    .searchSpace_0_write_data_din(in_36_write_data__din),
    .searchSpace_0_write_data_full_n(in_36_write_data__full_n),
    .searchSpace_0_write_data_write(in_36_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_36_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_36_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_36_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_36_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_36_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_36__din),
    .out_dist_full_n(out_dist_36__full_n),
    .out_dist_write(out_dist_36__write),
    .out_id_din(out_id_36__din),
    .out_id_full_n(out_id_36__full_n),
    .out_id_write(out_id_36__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_37
  krnl_partialKnn_wrapper_37_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_37_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_37_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_37_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_37_0__ap_ready),
    .start_id_0(64'd303104),
    .searchSpace_0_read_addr_s_din(in_37_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_37_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_37_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_37_0___in_37__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_37_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_37_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_37_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_37_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_37_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_37_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_37_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_37_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_37_0___in_37__q0),
    .searchSpace_0_write_data_din(in_37_write_data__din),
    .searchSpace_0_write_data_full_n(in_37_write_data__full_n),
    .searchSpace_0_write_data_write(in_37_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_37_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_37_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_37_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_37_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_37_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_37__din),
    .out_dist_full_n(out_dist_37__full_n),
    .out_dist_write(out_dist_37__write),
    .out_id_din(out_id_37__din),
    .out_id_full_n(out_id_37__full_n),
    .out_id_write(out_id_37__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_38
  krnl_partialKnn_wrapper_38_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_38_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_38_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_38_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_38_0__ap_ready),
    .start_id_0(64'd311296),
    .searchSpace_0_read_addr_s_din(in_38_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_38_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_38_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_38_0___in_38__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_38_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_38_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_38_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_38_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_38_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_38_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_38_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_38_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_38_0___in_38__q0),
    .searchSpace_0_write_data_din(in_38_write_data__din),
    .searchSpace_0_write_data_full_n(in_38_write_data__full_n),
    .searchSpace_0_write_data_write(in_38_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_38_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_38_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_38_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_38_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_38_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_38__din),
    .out_dist_full_n(out_dist_38__full_n),
    .out_dist_write(out_dist_38__write),
    .out_id_din(out_id_38__din),
    .out_id_full_n(out_id_38__full_n),
    .out_id_write(out_id_38__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_39
  krnl_partialKnn_wrapper_39_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_39_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_39_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_39_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_39_0__ap_ready),
    .start_id_0(64'd319488),
    .searchSpace_0_read_addr_s_din(in_39_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_39_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_39_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_39_0___in_39__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_39_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_39_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_39_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_39_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_39_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_39_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_39_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_39_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_39_0___in_39__q0),
    .searchSpace_0_write_data_din(in_39_write_data__din),
    .searchSpace_0_write_data_full_n(in_39_write_data__full_n),
    .searchSpace_0_write_data_write(in_39_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_39_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_39_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_39_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_39_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_39_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_39__din),
    .out_dist_full_n(out_dist_39__full_n),
    .out_dist_write(out_dist_39__write),
    .out_id_din(out_id_39__din),
    .out_id_full_n(out_id_39__full_n),
    .out_id_write(out_id_39__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_4
  krnl_partialKnn_wrapper_4_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_4_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_4_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_4_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_4_0__ap_ready),
    .start_id_0(64'd32768),
    .searchSpace_0_read_addr_s_din(in_4_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_4_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_4_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_4_0___in_4__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_4_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_4_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_4_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_4_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_4_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_4_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_4_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_4_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_4_0___in_4__q0),
    .searchSpace_0_write_data_din(in_4_write_data__din),
    .searchSpace_0_write_data_full_n(in_4_write_data__full_n),
    .searchSpace_0_write_data_write(in_4_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_4_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_4_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_4_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_4_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_4_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_4__din),
    .out_dist_full_n(out_dist_4__full_n),
    .out_dist_write(out_dist_4__write),
    .out_id_din(out_id_4__din),
    .out_id_full_n(out_id_4__full_n),
    .out_id_write(out_id_4__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_40
  krnl_partialKnn_wrapper_40_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_40_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_40_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_40_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_40_0__ap_ready),
    .start_id_0(64'd327680),
    .searchSpace_0_read_addr_s_din(in_40_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_40_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_40_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_40_0___in_40__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_40_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_40_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_40_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_40_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_40_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_40_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_40_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_40_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_40_0___in_40__q0),
    .searchSpace_0_write_data_din(in_40_write_data__din),
    .searchSpace_0_write_data_full_n(in_40_write_data__full_n),
    .searchSpace_0_write_data_write(in_40_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_40_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_40_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_40_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_40_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_40_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_40__din),
    .out_dist_full_n(out_dist_40__full_n),
    .out_dist_write(out_dist_40__write),
    .out_id_din(out_id_40__din),
    .out_id_full_n(out_id_40__full_n),
    .out_id_write(out_id_40__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_41
  krnl_partialKnn_wrapper_41_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_41_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_41_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_41_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_41_0__ap_ready),
    .start_id_0(64'd335872),
    .searchSpace_0_read_addr_s_din(in_41_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_41_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_41_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_41_0___in_41__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_41_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_41_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_41_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_41_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_41_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_41_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_41_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_41_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_41_0___in_41__q0),
    .searchSpace_0_write_data_din(in_41_write_data__din),
    .searchSpace_0_write_data_full_n(in_41_write_data__full_n),
    .searchSpace_0_write_data_write(in_41_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_41_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_41_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_41_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_41_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_41_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_41__din),
    .out_dist_full_n(out_dist_41__full_n),
    .out_dist_write(out_dist_41__write),
    .out_id_din(out_id_41__din),
    .out_id_full_n(out_id_41__full_n),
    .out_id_write(out_id_41__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_42
  krnl_partialKnn_wrapper_42_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_42_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_42_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_42_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_42_0__ap_ready),
    .start_id_0(64'd344064),
    .searchSpace_0_read_addr_s_din(in_42_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_42_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_42_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_42_0___in_42__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_42_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_42_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_42_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_42_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_42_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_42_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_42_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_42_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_42_0___in_42__q0),
    .searchSpace_0_write_data_din(in_42_write_data__din),
    .searchSpace_0_write_data_full_n(in_42_write_data__full_n),
    .searchSpace_0_write_data_write(in_42_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_42_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_42_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_42_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_42_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_42_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_42__din),
    .out_dist_full_n(out_dist_42__full_n),
    .out_dist_write(out_dist_42__write),
    .out_id_din(out_id_42__din),
    .out_id_full_n(out_id_42__full_n),
    .out_id_write(out_id_42__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_43
  krnl_partialKnn_wrapper_43_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_43_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_43_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_43_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_43_0__ap_ready),
    .start_id_0(64'd352256),
    .searchSpace_0_read_addr_s_din(in_43_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_43_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_43_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_43_0___in_43__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_43_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_43_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_43_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_43_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_43_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_43_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_43_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_43_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_43_0___in_43__q0),
    .searchSpace_0_write_data_din(in_43_write_data__din),
    .searchSpace_0_write_data_full_n(in_43_write_data__full_n),
    .searchSpace_0_write_data_write(in_43_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_43_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_43_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_43_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_43_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_43_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_43__din),
    .out_dist_full_n(out_dist_43__full_n),
    .out_dist_write(out_dist_43__write),
    .out_id_din(out_id_43__din),
    .out_id_full_n(out_id_43__full_n),
    .out_id_write(out_id_43__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_44
  krnl_partialKnn_wrapper_44_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_44_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_44_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_44_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_44_0__ap_ready),
    .start_id_0(64'd360448),
    .searchSpace_0_read_addr_s_din(in_44_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_44_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_44_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_44_0___in_44__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_44_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_44_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_44_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_44_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_44_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_44_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_44_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_44_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_44_0___in_44__q0),
    .searchSpace_0_write_data_din(in_44_write_data__din),
    .searchSpace_0_write_data_full_n(in_44_write_data__full_n),
    .searchSpace_0_write_data_write(in_44_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_44_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_44_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_44_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_44_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_44_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_44__din),
    .out_dist_full_n(out_dist_44__full_n),
    .out_dist_write(out_dist_44__write),
    .out_id_din(out_id_44__din),
    .out_id_full_n(out_id_44__full_n),
    .out_id_write(out_id_44__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_45
  krnl_partialKnn_wrapper_45_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_45_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_45_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_45_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_45_0__ap_ready),
    .start_id_0(64'd368640),
    .searchSpace_0_read_addr_s_din(in_45_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_45_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_45_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_45_0___in_45__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_45_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_45_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_45_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_45_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_45_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_45_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_45_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_45_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_45_0___in_45__q0),
    .searchSpace_0_write_data_din(in_45_write_data__din),
    .searchSpace_0_write_data_full_n(in_45_write_data__full_n),
    .searchSpace_0_write_data_write(in_45_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_45_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_45_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_45_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_45_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_45_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_45__din),
    .out_dist_full_n(out_dist_45__full_n),
    .out_dist_write(out_dist_45__write),
    .out_id_din(out_id_45__din),
    .out_id_full_n(out_id_45__full_n),
    .out_id_write(out_id_45__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_46
  krnl_partialKnn_wrapper_46_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_46_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_46_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_46_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_46_0__ap_ready),
    .start_id_0(64'd376832),
    .searchSpace_0_read_addr_s_din(in_46_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_46_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_46_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_46_0___in_46__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_46_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_46_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_46_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_46_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_46_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_46_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_46_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_46_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_46_0___in_46__q0),
    .searchSpace_0_write_data_din(in_46_write_data__din),
    .searchSpace_0_write_data_full_n(in_46_write_data__full_n),
    .searchSpace_0_write_data_write(in_46_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_46_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_46_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_46_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_46_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_46_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_46__din),
    .out_dist_full_n(out_dist_46__full_n),
    .out_dist_write(out_dist_46__write),
    .out_id_din(out_id_46__din),
    .out_id_full_n(out_id_46__full_n),
    .out_id_write(out_id_46__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_47
  krnl_partialKnn_wrapper_47_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_47_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_47_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_47_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_47_0__ap_ready),
    .start_id_0(64'd385024),
    .searchSpace_0_read_addr_s_din(in_47_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_47_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_47_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_47_0___in_47__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_47_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_47_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_47_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_47_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_47_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_47_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_47_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_47_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_47_0___in_47__q0),
    .searchSpace_0_write_data_din(in_47_write_data__din),
    .searchSpace_0_write_data_full_n(in_47_write_data__full_n),
    .searchSpace_0_write_data_write(in_47_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_47_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_47_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_47_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_47_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_47_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_47__din),
    .out_dist_full_n(out_dist_47__full_n),
    .out_dist_write(out_dist_47__write),
    .out_id_din(out_id_47__din),
    .out_id_full_n(out_id_47__full_n),
    .out_id_write(out_id_47__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_48
  krnl_partialKnn_wrapper_48_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_48_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_48_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_48_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_48_0__ap_ready),
    .start_id_0(64'd393216),
    .searchSpace_0_read_addr_s_din(in_48_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_48_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_48_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_48_0___in_48__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_48_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_48_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_48_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_48_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_48_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_48_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_48_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_48_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_48_0___in_48__q0),
    .searchSpace_0_write_data_din(in_48_write_data__din),
    .searchSpace_0_write_data_full_n(in_48_write_data__full_n),
    .searchSpace_0_write_data_write(in_48_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_48_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_48_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_48_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_48_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_48_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_48__din),
    .out_dist_full_n(out_dist_48__full_n),
    .out_dist_write(out_dist_48__write),
    .out_id_din(out_id_48__din),
    .out_id_full_n(out_id_48__full_n),
    .out_id_write(out_id_48__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_49
  krnl_partialKnn_wrapper_49_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_49_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_49_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_49_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_49_0__ap_ready),
    .start_id_0(64'd401408),
    .searchSpace_0_read_addr_s_din(in_49_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_49_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_49_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_49_0___in_49__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_49_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_49_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_49_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_49_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_49_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_49_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_49_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_49_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_49_0___in_49__q0),
    .searchSpace_0_write_data_din(in_49_write_data__din),
    .searchSpace_0_write_data_full_n(in_49_write_data__full_n),
    .searchSpace_0_write_data_write(in_49_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_49_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_49_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_49_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_49_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_49_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_49__din),
    .out_dist_full_n(out_dist_49__full_n),
    .out_dist_write(out_dist_49__write),
    .out_id_din(out_id_49__din),
    .out_id_full_n(out_id_49__full_n),
    .out_id_write(out_id_49__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_5
  krnl_partialKnn_wrapper_5_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_5_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_5_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_5_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_5_0__ap_ready),
    .start_id_0(64'd40960),
    .searchSpace_0_read_addr_s_din(in_5_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_5_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_5_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_5_0___in_5__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_5_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_5_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_5_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_5_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_5_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_5_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_5_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_5_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_5_0___in_5__q0),
    .searchSpace_0_write_data_din(in_5_write_data__din),
    .searchSpace_0_write_data_full_n(in_5_write_data__full_n),
    .searchSpace_0_write_data_write(in_5_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_5_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_5_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_5_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_5_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_5_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_5__din),
    .out_dist_full_n(out_dist_5__full_n),
    .out_dist_write(out_dist_5__write),
    .out_id_din(out_id_5__din),
    .out_id_full_n(out_id_5__full_n),
    .out_id_write(out_id_5__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_50
  krnl_partialKnn_wrapper_50_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_50_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_50_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_50_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_50_0__ap_ready),
    .start_id_0(64'd409600),
    .searchSpace_0_read_addr_s_din(in_50_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_50_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_50_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_50_0___in_50__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_50_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_50_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_50_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_50_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_50_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_50_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_50_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_50_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_50_0___in_50__q0),
    .searchSpace_0_write_data_din(in_50_write_data__din),
    .searchSpace_0_write_data_full_n(in_50_write_data__full_n),
    .searchSpace_0_write_data_write(in_50_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_50_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_50_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_50_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_50_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_50_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_50__din),
    .out_dist_full_n(out_dist_50__full_n),
    .out_dist_write(out_dist_50__write),
    .out_id_din(out_id_50__din),
    .out_id_full_n(out_id_50__full_n),
    .out_id_write(out_id_50__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_51
  krnl_partialKnn_wrapper_51_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_51_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_51_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_51_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_51_0__ap_ready),
    .start_id_0(64'd417792),
    .searchSpace_0_read_addr_s_din(in_51_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_51_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_51_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_51_0___in_51__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_51_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_51_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_51_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_51_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_51_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_51_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_51_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_51_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_51_0___in_51__q0),
    .searchSpace_0_write_data_din(in_51_write_data__din),
    .searchSpace_0_write_data_full_n(in_51_write_data__full_n),
    .searchSpace_0_write_data_write(in_51_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_51_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_51_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_51_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_51_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_51_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_51__din),
    .out_dist_full_n(out_dist_51__full_n),
    .out_dist_write(out_dist_51__write),
    .out_id_din(out_id_51__din),
    .out_id_full_n(out_id_51__full_n),
    .out_id_write(out_id_51__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_52
  krnl_partialKnn_wrapper_52_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_52_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_52_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_52_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_52_0__ap_ready),
    .start_id_0(64'd425984),
    .searchSpace_0_read_addr_s_din(in_52_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_52_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_52_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_52_0___in_52__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_52_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_52_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_52_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_52_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_52_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_52_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_52_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_52_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_52_0___in_52__q0),
    .searchSpace_0_write_data_din(in_52_write_data__din),
    .searchSpace_0_write_data_full_n(in_52_write_data__full_n),
    .searchSpace_0_write_data_write(in_52_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_52_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_52_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_52_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_52_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_52_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_52__din),
    .out_dist_full_n(out_dist_52__full_n),
    .out_dist_write(out_dist_52__write),
    .out_id_din(out_id_52__din),
    .out_id_full_n(out_id_52__full_n),
    .out_id_write(out_id_52__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_53
  krnl_partialKnn_wrapper_53_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_53_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_53_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_53_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_53_0__ap_ready),
    .start_id_0(64'd434176),
    .searchSpace_0_read_addr_s_din(in_53_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_53_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_53_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_53_0___in_53__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_53_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_53_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_53_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_53_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_53_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_53_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_53_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_53_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_53_0___in_53__q0),
    .searchSpace_0_write_data_din(in_53_write_data__din),
    .searchSpace_0_write_data_full_n(in_53_write_data__full_n),
    .searchSpace_0_write_data_write(in_53_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_53_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_53_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_53_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_53_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_53_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_53__din),
    .out_dist_full_n(out_dist_53__full_n),
    .out_dist_write(out_dist_53__write),
    .out_id_din(out_id_53__din),
    .out_id_full_n(out_id_53__full_n),
    .out_id_write(out_id_53__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_6
  krnl_partialKnn_wrapper_6_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_6_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_6_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_6_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_6_0__ap_ready),
    .start_id_0(64'd49152),
    .searchSpace_0_read_addr_s_din(in_6_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_6_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_6_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_6_0___in_6__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_6_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_6_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_6_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_6_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_6_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_6_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_6_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_6_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_6_0___in_6__q0),
    .searchSpace_0_write_data_din(in_6_write_data__din),
    .searchSpace_0_write_data_full_n(in_6_write_data__full_n),
    .searchSpace_0_write_data_write(in_6_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_6_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_6_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_6_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_6_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_6_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_6__din),
    .out_dist_full_n(out_dist_6__full_n),
    .out_dist_write(out_dist_6__write),
    .out_id_din(out_id_6__din),
    .out_id_full_n(out_id_6__full_n),
    .out_id_write(out_id_6__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_7
  krnl_partialKnn_wrapper_7_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_7_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_7_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_7_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_7_0__ap_ready),
    .start_id_0(64'd57344),
    .searchSpace_0_read_addr_s_din(in_7_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_7_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_7_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_7_0___in_7__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_7_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_7_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_7_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_7_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_7_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_7_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_7_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_7_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_7_0___in_7__q0),
    .searchSpace_0_write_data_din(in_7_write_data__din),
    .searchSpace_0_write_data_full_n(in_7_write_data__full_n),
    .searchSpace_0_write_data_write(in_7_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_7_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_7_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_7_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_7_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_7_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_7__din),
    .out_dist_full_n(out_dist_7__full_n),
    .out_dist_write(out_dist_7__write),
    .out_id_din(out_id_7__din),
    .out_id_full_n(out_id_7__full_n),
    .out_id_write(out_id_7__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_8
  krnl_partialKnn_wrapper_8_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_8_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_8_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_8_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_8_0__ap_ready),
    .start_id_0(64'd65536),
    .searchSpace_0_read_addr_s_din(in_8_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_8_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_8_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_8_0___in_8__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_8_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_8_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_8_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_8_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_8_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_8_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_8_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_8_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_8_0___in_8__q0),
    .searchSpace_0_write_data_din(in_8_write_data__din),
    .searchSpace_0_write_data_full_n(in_8_write_data__full_n),
    .searchSpace_0_write_data_write(in_8_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_8_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_8_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_8_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_8_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_8_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_8__din),
    .out_dist_full_n(out_dist_8__full_n),
    .out_dist_write(out_dist_8__write),
    .out_id_din(out_id_8__din),
    .out_id_full_n(out_id_8__full_n),
    .out_id_write(out_id_8__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_9
  krnl_partialKnn_wrapper_9_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_9_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_9_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_9_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_9_0__ap_ready),
    .start_id_0(64'd73728),
    .searchSpace_0_read_addr_s_din(in_9_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_9_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_9_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_9_0___in_9__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_9_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_9_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_9_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_9_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_9_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_9_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_9_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_9_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_9_0___in_9__q0),
    .searchSpace_0_write_data_din(in_9_write_data__din),
    .searchSpace_0_write_data_full_n(in_9_write_data__full_n),
    .searchSpace_0_write_data_write(in_9_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_9_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_9_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_9_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_9_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_9_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_9__din),
    .out_dist_full_n(out_dist_9__full_n),
    .out_dist_write(out_dist_9__write),
    .out_id_din(out_id_9__din),
    .out_id_full_n(out_id_9__full_n),
    .out_id_write(out_id_9__write)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(32),
    .DataWidthBytesLog(2),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(255)
  )
  L4_out_dist__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_L4_out_dist_ARADDR),
    .m_axi_ARBURST(m_axi_L4_out_dist_ARBURST),
    .m_axi_ARCACHE(m_axi_L4_out_dist_ARCACHE),
    .m_axi_ARID(m_axi_L4_out_dist_ARID),
    .m_axi_ARLEN(m_axi_L4_out_dist_ARLEN),
    .m_axi_ARLOCK(m_axi_L4_out_dist_ARLOCK),
    .m_axi_ARPROT(m_axi_L4_out_dist_ARPROT),
    .m_axi_ARQOS(m_axi_L4_out_dist_ARQOS),
    .m_axi_ARREADY(m_axi_L4_out_dist_ARREADY),
    .m_axi_ARSIZE(m_axi_L4_out_dist_ARSIZE),
    .m_axi_ARVALID(m_axi_L4_out_dist_ARVALID),
    .m_axi_AWADDR(m_axi_L4_out_dist_AWADDR),
    .m_axi_AWBURST(m_axi_L4_out_dist_AWBURST),
    .m_axi_AWCACHE(m_axi_L4_out_dist_AWCACHE),
    .m_axi_AWID(m_axi_L4_out_dist_AWID),
    .m_axi_AWLEN(m_axi_L4_out_dist_AWLEN),
    .m_axi_AWLOCK(m_axi_L4_out_dist_AWLOCK),
    .m_axi_AWPROT(m_axi_L4_out_dist_AWPROT),
    .m_axi_AWQOS(m_axi_L4_out_dist_AWQOS),
    .m_axi_AWREADY(m_axi_L4_out_dist_AWREADY),
    .m_axi_AWSIZE(m_axi_L4_out_dist_AWSIZE),
    .m_axi_AWVALID(m_axi_L4_out_dist_AWVALID),
    .m_axi_BID(m_axi_L4_out_dist_BID),
    .m_axi_BREADY(m_axi_L4_out_dist_BREADY),
    .m_axi_BRESP(m_axi_L4_out_dist_BRESP),
    .m_axi_BVALID(m_axi_L4_out_dist_BVALID),
    .m_axi_RDATA(m_axi_L4_out_dist_RDATA),
    .m_axi_RID(m_axi_L4_out_dist_RID),
    .m_axi_RLAST(m_axi_L4_out_dist_RLAST),
    .m_axi_RREADY(m_axi_L4_out_dist_RREADY),
    .m_axi_RRESP(m_axi_L4_out_dist_RRESP),
    .m_axi_RVALID(m_axi_L4_out_dist_RVALID),
    .m_axi_WDATA(m_axi_L4_out_dist_WDATA),
    .m_axi_WLAST(m_axi_L4_out_dist_WLAST),
    .m_axi_WREADY(m_axi_L4_out_dist_WREADY),
    .m_axi_WSTRB(m_axi_L4_out_dist_WSTRB),
    .m_axi_WVALID(m_axi_L4_out_dist_WVALID),
    .read_addr_din(L4_out_dist_read_addr__din),
    .read_addr_full_n(L4_out_dist_read_addr__full_n),
    .read_addr_write(L4_out_dist_read_addr__write),
    .read_data_dout(L4_out_dist_read_data__dout),
    .read_data_empty_n(L4_out_dist_read_data__empty_n),
    .read_data_read(L4_out_dist_read_data__read),
    .write_addr_din(L4_out_dist_write_addr__din),
    .write_addr_full_n(L4_out_dist_write_addr__full_n),
    .write_addr_write(L4_out_dist_write_addr__write),
    .write_data_din(L4_out_dist_write_data__din),
    .write_data_full_n(L4_out_dist_write_data__full_n),
    .write_data_write(L4_out_dist_write_data__write),
    .write_resp_dout(L4_out_dist_write_resp__dout),
    .write_resp_empty_n(L4_out_dist_write_resp__empty_n),
    .write_resp_read(L4_out_dist_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(32),
    .DataWidthBytesLog(2),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(255)
  )
  L4_out_id__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_L4_out_id_ARADDR),
    .m_axi_ARBURST(m_axi_L4_out_id_ARBURST),
    .m_axi_ARCACHE(m_axi_L4_out_id_ARCACHE),
    .m_axi_ARID(m_axi_L4_out_id_ARID),
    .m_axi_ARLEN(m_axi_L4_out_id_ARLEN),
    .m_axi_ARLOCK(m_axi_L4_out_id_ARLOCK),
    .m_axi_ARPROT(m_axi_L4_out_id_ARPROT),
    .m_axi_ARQOS(m_axi_L4_out_id_ARQOS),
    .m_axi_ARREADY(m_axi_L4_out_id_ARREADY),
    .m_axi_ARSIZE(m_axi_L4_out_id_ARSIZE),
    .m_axi_ARVALID(m_axi_L4_out_id_ARVALID),
    .m_axi_AWADDR(m_axi_L4_out_id_AWADDR),
    .m_axi_AWBURST(m_axi_L4_out_id_AWBURST),
    .m_axi_AWCACHE(m_axi_L4_out_id_AWCACHE),
    .m_axi_AWID(m_axi_L4_out_id_AWID),
    .m_axi_AWLEN(m_axi_L4_out_id_AWLEN),
    .m_axi_AWLOCK(m_axi_L4_out_id_AWLOCK),
    .m_axi_AWPROT(m_axi_L4_out_id_AWPROT),
    .m_axi_AWQOS(m_axi_L4_out_id_AWQOS),
    .m_axi_AWREADY(m_axi_L4_out_id_AWREADY),
    .m_axi_AWSIZE(m_axi_L4_out_id_AWSIZE),
    .m_axi_AWVALID(m_axi_L4_out_id_AWVALID),
    .m_axi_BID(m_axi_L4_out_id_BID),
    .m_axi_BREADY(m_axi_L4_out_id_BREADY),
    .m_axi_BRESP(m_axi_L4_out_id_BRESP),
    .m_axi_BVALID(m_axi_L4_out_id_BVALID),
    .m_axi_RDATA(m_axi_L4_out_id_RDATA),
    .m_axi_RID(m_axi_L4_out_id_RID),
    .m_axi_RLAST(m_axi_L4_out_id_RLAST),
    .m_axi_RREADY(m_axi_L4_out_id_RREADY),
    .m_axi_RRESP(m_axi_L4_out_id_RRESP),
    .m_axi_RVALID(m_axi_L4_out_id_RVALID),
    .m_axi_WDATA(m_axi_L4_out_id_WDATA),
    .m_axi_WLAST(m_axi_L4_out_id_WLAST),
    .m_axi_WREADY(m_axi_L4_out_id_WREADY),
    .m_axi_WSTRB(m_axi_L4_out_id_WSTRB),
    .m_axi_WVALID(m_axi_L4_out_id_WVALID),
    .read_addr_din(L4_out_id_read_addr__din),
    .read_addr_full_n(L4_out_id_read_addr__full_n),
    .read_addr_write(L4_out_id_read_addr__write),
    .read_data_dout(L4_out_id_read_data__dout),
    .read_data_empty_n(L4_out_id_read_data__empty_n),
    .read_data_read(L4_out_id_read_data__read),
    .write_addr_din(L4_out_id_write_addr__din),
    .write_addr_full_n(L4_out_id_write_addr__full_n),
    .write_addr_write(L4_out_id_write_addr__write),
    .write_data_din(L4_out_id_write_data__din),
    .write_data_full_n(L4_out_id_write_data__full_n),
    .write_data_write(L4_out_id_write_data__write),
    .write_resp_dout(L4_out_id_write_resp__dout),
    .write_resp_empty_n(L4_out_id_write_resp__empty_n),
    .write_resp_read(L4_out_id_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_0_ARADDR),
    .m_axi_ARBURST(m_axi_in_0_ARBURST),
    .m_axi_ARCACHE(m_axi_in_0_ARCACHE),
    .m_axi_ARID(m_axi_in_0_ARID),
    .m_axi_ARLEN(m_axi_in_0_ARLEN),
    .m_axi_ARLOCK(m_axi_in_0_ARLOCK),
    .m_axi_ARPROT(m_axi_in_0_ARPROT),
    .m_axi_ARQOS(m_axi_in_0_ARQOS),
    .m_axi_ARREADY(m_axi_in_0_ARREADY),
    .m_axi_ARSIZE(m_axi_in_0_ARSIZE),
    .m_axi_ARVALID(m_axi_in_0_ARVALID),
    .m_axi_AWADDR(m_axi_in_0_AWADDR),
    .m_axi_AWBURST(m_axi_in_0_AWBURST),
    .m_axi_AWCACHE(m_axi_in_0_AWCACHE),
    .m_axi_AWID(m_axi_in_0_AWID),
    .m_axi_AWLEN(m_axi_in_0_AWLEN),
    .m_axi_AWLOCK(m_axi_in_0_AWLOCK),
    .m_axi_AWPROT(m_axi_in_0_AWPROT),
    .m_axi_AWQOS(m_axi_in_0_AWQOS),
    .m_axi_AWREADY(m_axi_in_0_AWREADY),
    .m_axi_AWSIZE(m_axi_in_0_AWSIZE),
    .m_axi_AWVALID(m_axi_in_0_AWVALID),
    .m_axi_BID(m_axi_in_0_BID),
    .m_axi_BREADY(m_axi_in_0_BREADY),
    .m_axi_BRESP(m_axi_in_0_BRESP),
    .m_axi_BVALID(m_axi_in_0_BVALID),
    .m_axi_RDATA(m_axi_in_0_RDATA),
    .m_axi_RID(m_axi_in_0_RID),
    .m_axi_RLAST(m_axi_in_0_RLAST),
    .m_axi_RREADY(m_axi_in_0_RREADY),
    .m_axi_RRESP(m_axi_in_0_RRESP),
    .m_axi_RVALID(m_axi_in_0_RVALID),
    .m_axi_WDATA(m_axi_in_0_WDATA),
    .m_axi_WLAST(m_axi_in_0_WLAST),
    .m_axi_WREADY(m_axi_in_0_WREADY),
    .m_axi_WSTRB(m_axi_in_0_WSTRB),
    .m_axi_WVALID(m_axi_in_0_WVALID),
    .read_addr_din(in_0_read_addr__din),
    .read_addr_full_n(in_0_read_addr__full_n),
    .read_addr_write(in_0_read_addr__write),
    .read_data_dout(in_0_read_data__dout),
    .read_data_empty_n(in_0_read_data__empty_n),
    .read_data_read(in_0_read_data__read),
    .write_addr_din(in_0_write_addr__din),
    .write_addr_full_n(in_0_write_addr__full_n),
    .write_addr_write(in_0_write_addr__write),
    .write_data_din(in_0_write_data__din),
    .write_data_full_n(in_0_write_data__full_n),
    .write_data_write(in_0_write_data__write),
    .write_resp_dout(in_0_write_resp__dout),
    .write_resp_empty_n(in_0_write_resp__empty_n),
    .write_resp_read(in_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_1_ARADDR),
    .m_axi_ARBURST(m_axi_in_1_ARBURST),
    .m_axi_ARCACHE(m_axi_in_1_ARCACHE),
    .m_axi_ARID(m_axi_in_1_ARID),
    .m_axi_ARLEN(m_axi_in_1_ARLEN),
    .m_axi_ARLOCK(m_axi_in_1_ARLOCK),
    .m_axi_ARPROT(m_axi_in_1_ARPROT),
    .m_axi_ARQOS(m_axi_in_1_ARQOS),
    .m_axi_ARREADY(m_axi_in_1_ARREADY),
    .m_axi_ARSIZE(m_axi_in_1_ARSIZE),
    .m_axi_ARVALID(m_axi_in_1_ARVALID),
    .m_axi_AWADDR(m_axi_in_1_AWADDR),
    .m_axi_AWBURST(m_axi_in_1_AWBURST),
    .m_axi_AWCACHE(m_axi_in_1_AWCACHE),
    .m_axi_AWID(m_axi_in_1_AWID),
    .m_axi_AWLEN(m_axi_in_1_AWLEN),
    .m_axi_AWLOCK(m_axi_in_1_AWLOCK),
    .m_axi_AWPROT(m_axi_in_1_AWPROT),
    .m_axi_AWQOS(m_axi_in_1_AWQOS),
    .m_axi_AWREADY(m_axi_in_1_AWREADY),
    .m_axi_AWSIZE(m_axi_in_1_AWSIZE),
    .m_axi_AWVALID(m_axi_in_1_AWVALID),
    .m_axi_BID(m_axi_in_1_BID),
    .m_axi_BREADY(m_axi_in_1_BREADY),
    .m_axi_BRESP(m_axi_in_1_BRESP),
    .m_axi_BVALID(m_axi_in_1_BVALID),
    .m_axi_RDATA(m_axi_in_1_RDATA),
    .m_axi_RID(m_axi_in_1_RID),
    .m_axi_RLAST(m_axi_in_1_RLAST),
    .m_axi_RREADY(m_axi_in_1_RREADY),
    .m_axi_RRESP(m_axi_in_1_RRESP),
    .m_axi_RVALID(m_axi_in_1_RVALID),
    .m_axi_WDATA(m_axi_in_1_WDATA),
    .m_axi_WLAST(m_axi_in_1_WLAST),
    .m_axi_WREADY(m_axi_in_1_WREADY),
    .m_axi_WSTRB(m_axi_in_1_WSTRB),
    .m_axi_WVALID(m_axi_in_1_WVALID),
    .read_addr_din(in_1_read_addr__din),
    .read_addr_full_n(in_1_read_addr__full_n),
    .read_addr_write(in_1_read_addr__write),
    .read_data_dout(in_1_read_data__dout),
    .read_data_empty_n(in_1_read_data__empty_n),
    .read_data_read(in_1_read_data__read),
    .write_addr_din(in_1_write_addr__din),
    .write_addr_full_n(in_1_write_addr__full_n),
    .write_addr_write(in_1_write_addr__write),
    .write_data_din(in_1_write_data__din),
    .write_data_full_n(in_1_write_data__full_n),
    .write_data_write(in_1_write_data__write),
    .write_resp_dout(in_1_write_resp__dout),
    .write_resp_empty_n(in_1_write_resp__empty_n),
    .write_resp_read(in_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_10__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_10_ARADDR),
    .m_axi_ARBURST(m_axi_in_10_ARBURST),
    .m_axi_ARCACHE(m_axi_in_10_ARCACHE),
    .m_axi_ARID(m_axi_in_10_ARID),
    .m_axi_ARLEN(m_axi_in_10_ARLEN),
    .m_axi_ARLOCK(m_axi_in_10_ARLOCK),
    .m_axi_ARPROT(m_axi_in_10_ARPROT),
    .m_axi_ARQOS(m_axi_in_10_ARQOS),
    .m_axi_ARREADY(m_axi_in_10_ARREADY),
    .m_axi_ARSIZE(m_axi_in_10_ARSIZE),
    .m_axi_ARVALID(m_axi_in_10_ARVALID),
    .m_axi_AWADDR(m_axi_in_10_AWADDR),
    .m_axi_AWBURST(m_axi_in_10_AWBURST),
    .m_axi_AWCACHE(m_axi_in_10_AWCACHE),
    .m_axi_AWID(m_axi_in_10_AWID),
    .m_axi_AWLEN(m_axi_in_10_AWLEN),
    .m_axi_AWLOCK(m_axi_in_10_AWLOCK),
    .m_axi_AWPROT(m_axi_in_10_AWPROT),
    .m_axi_AWQOS(m_axi_in_10_AWQOS),
    .m_axi_AWREADY(m_axi_in_10_AWREADY),
    .m_axi_AWSIZE(m_axi_in_10_AWSIZE),
    .m_axi_AWVALID(m_axi_in_10_AWVALID),
    .m_axi_BID(m_axi_in_10_BID),
    .m_axi_BREADY(m_axi_in_10_BREADY),
    .m_axi_BRESP(m_axi_in_10_BRESP),
    .m_axi_BVALID(m_axi_in_10_BVALID),
    .m_axi_RDATA(m_axi_in_10_RDATA),
    .m_axi_RID(m_axi_in_10_RID),
    .m_axi_RLAST(m_axi_in_10_RLAST),
    .m_axi_RREADY(m_axi_in_10_RREADY),
    .m_axi_RRESP(m_axi_in_10_RRESP),
    .m_axi_RVALID(m_axi_in_10_RVALID),
    .m_axi_WDATA(m_axi_in_10_WDATA),
    .m_axi_WLAST(m_axi_in_10_WLAST),
    .m_axi_WREADY(m_axi_in_10_WREADY),
    .m_axi_WSTRB(m_axi_in_10_WSTRB),
    .m_axi_WVALID(m_axi_in_10_WVALID),
    .read_addr_din(in_10_read_addr__din),
    .read_addr_full_n(in_10_read_addr__full_n),
    .read_addr_write(in_10_read_addr__write),
    .read_data_dout(in_10_read_data__dout),
    .read_data_empty_n(in_10_read_data__empty_n),
    .read_data_read(in_10_read_data__read),
    .write_addr_din(in_10_write_addr__din),
    .write_addr_full_n(in_10_write_addr__full_n),
    .write_addr_write(in_10_write_addr__write),
    .write_data_din(in_10_write_data__din),
    .write_data_full_n(in_10_write_data__full_n),
    .write_data_write(in_10_write_data__write),
    .write_resp_dout(in_10_write_resp__dout),
    .write_resp_empty_n(in_10_write_resp__empty_n),
    .write_resp_read(in_10_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_11__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_11_ARADDR),
    .m_axi_ARBURST(m_axi_in_11_ARBURST),
    .m_axi_ARCACHE(m_axi_in_11_ARCACHE),
    .m_axi_ARID(m_axi_in_11_ARID),
    .m_axi_ARLEN(m_axi_in_11_ARLEN),
    .m_axi_ARLOCK(m_axi_in_11_ARLOCK),
    .m_axi_ARPROT(m_axi_in_11_ARPROT),
    .m_axi_ARQOS(m_axi_in_11_ARQOS),
    .m_axi_ARREADY(m_axi_in_11_ARREADY),
    .m_axi_ARSIZE(m_axi_in_11_ARSIZE),
    .m_axi_ARVALID(m_axi_in_11_ARVALID),
    .m_axi_AWADDR(m_axi_in_11_AWADDR),
    .m_axi_AWBURST(m_axi_in_11_AWBURST),
    .m_axi_AWCACHE(m_axi_in_11_AWCACHE),
    .m_axi_AWID(m_axi_in_11_AWID),
    .m_axi_AWLEN(m_axi_in_11_AWLEN),
    .m_axi_AWLOCK(m_axi_in_11_AWLOCK),
    .m_axi_AWPROT(m_axi_in_11_AWPROT),
    .m_axi_AWQOS(m_axi_in_11_AWQOS),
    .m_axi_AWREADY(m_axi_in_11_AWREADY),
    .m_axi_AWSIZE(m_axi_in_11_AWSIZE),
    .m_axi_AWVALID(m_axi_in_11_AWVALID),
    .m_axi_BID(m_axi_in_11_BID),
    .m_axi_BREADY(m_axi_in_11_BREADY),
    .m_axi_BRESP(m_axi_in_11_BRESP),
    .m_axi_BVALID(m_axi_in_11_BVALID),
    .m_axi_RDATA(m_axi_in_11_RDATA),
    .m_axi_RID(m_axi_in_11_RID),
    .m_axi_RLAST(m_axi_in_11_RLAST),
    .m_axi_RREADY(m_axi_in_11_RREADY),
    .m_axi_RRESP(m_axi_in_11_RRESP),
    .m_axi_RVALID(m_axi_in_11_RVALID),
    .m_axi_WDATA(m_axi_in_11_WDATA),
    .m_axi_WLAST(m_axi_in_11_WLAST),
    .m_axi_WREADY(m_axi_in_11_WREADY),
    .m_axi_WSTRB(m_axi_in_11_WSTRB),
    .m_axi_WVALID(m_axi_in_11_WVALID),
    .read_addr_din(in_11_read_addr__din),
    .read_addr_full_n(in_11_read_addr__full_n),
    .read_addr_write(in_11_read_addr__write),
    .read_data_dout(in_11_read_data__dout),
    .read_data_empty_n(in_11_read_data__empty_n),
    .read_data_read(in_11_read_data__read),
    .write_addr_din(in_11_write_addr__din),
    .write_addr_full_n(in_11_write_addr__full_n),
    .write_addr_write(in_11_write_addr__write),
    .write_data_din(in_11_write_data__din),
    .write_data_full_n(in_11_write_data__full_n),
    .write_data_write(in_11_write_data__write),
    .write_resp_dout(in_11_write_resp__dout),
    .write_resp_empty_n(in_11_write_resp__empty_n),
    .write_resp_read(in_11_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_12__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_12_ARADDR),
    .m_axi_ARBURST(m_axi_in_12_ARBURST),
    .m_axi_ARCACHE(m_axi_in_12_ARCACHE),
    .m_axi_ARID(m_axi_in_12_ARID),
    .m_axi_ARLEN(m_axi_in_12_ARLEN),
    .m_axi_ARLOCK(m_axi_in_12_ARLOCK),
    .m_axi_ARPROT(m_axi_in_12_ARPROT),
    .m_axi_ARQOS(m_axi_in_12_ARQOS),
    .m_axi_ARREADY(m_axi_in_12_ARREADY),
    .m_axi_ARSIZE(m_axi_in_12_ARSIZE),
    .m_axi_ARVALID(m_axi_in_12_ARVALID),
    .m_axi_AWADDR(m_axi_in_12_AWADDR),
    .m_axi_AWBURST(m_axi_in_12_AWBURST),
    .m_axi_AWCACHE(m_axi_in_12_AWCACHE),
    .m_axi_AWID(m_axi_in_12_AWID),
    .m_axi_AWLEN(m_axi_in_12_AWLEN),
    .m_axi_AWLOCK(m_axi_in_12_AWLOCK),
    .m_axi_AWPROT(m_axi_in_12_AWPROT),
    .m_axi_AWQOS(m_axi_in_12_AWQOS),
    .m_axi_AWREADY(m_axi_in_12_AWREADY),
    .m_axi_AWSIZE(m_axi_in_12_AWSIZE),
    .m_axi_AWVALID(m_axi_in_12_AWVALID),
    .m_axi_BID(m_axi_in_12_BID),
    .m_axi_BREADY(m_axi_in_12_BREADY),
    .m_axi_BRESP(m_axi_in_12_BRESP),
    .m_axi_BVALID(m_axi_in_12_BVALID),
    .m_axi_RDATA(m_axi_in_12_RDATA),
    .m_axi_RID(m_axi_in_12_RID),
    .m_axi_RLAST(m_axi_in_12_RLAST),
    .m_axi_RREADY(m_axi_in_12_RREADY),
    .m_axi_RRESP(m_axi_in_12_RRESP),
    .m_axi_RVALID(m_axi_in_12_RVALID),
    .m_axi_WDATA(m_axi_in_12_WDATA),
    .m_axi_WLAST(m_axi_in_12_WLAST),
    .m_axi_WREADY(m_axi_in_12_WREADY),
    .m_axi_WSTRB(m_axi_in_12_WSTRB),
    .m_axi_WVALID(m_axi_in_12_WVALID),
    .read_addr_din(in_12_read_addr__din),
    .read_addr_full_n(in_12_read_addr__full_n),
    .read_addr_write(in_12_read_addr__write),
    .read_data_dout(in_12_read_data__dout),
    .read_data_empty_n(in_12_read_data__empty_n),
    .read_data_read(in_12_read_data__read),
    .write_addr_din(in_12_write_addr__din),
    .write_addr_full_n(in_12_write_addr__full_n),
    .write_addr_write(in_12_write_addr__write),
    .write_data_din(in_12_write_data__din),
    .write_data_full_n(in_12_write_data__full_n),
    .write_data_write(in_12_write_data__write),
    .write_resp_dout(in_12_write_resp__dout),
    .write_resp_empty_n(in_12_write_resp__empty_n),
    .write_resp_read(in_12_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_13__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_13_ARADDR),
    .m_axi_ARBURST(m_axi_in_13_ARBURST),
    .m_axi_ARCACHE(m_axi_in_13_ARCACHE),
    .m_axi_ARID(m_axi_in_13_ARID),
    .m_axi_ARLEN(m_axi_in_13_ARLEN),
    .m_axi_ARLOCK(m_axi_in_13_ARLOCK),
    .m_axi_ARPROT(m_axi_in_13_ARPROT),
    .m_axi_ARQOS(m_axi_in_13_ARQOS),
    .m_axi_ARREADY(m_axi_in_13_ARREADY),
    .m_axi_ARSIZE(m_axi_in_13_ARSIZE),
    .m_axi_ARVALID(m_axi_in_13_ARVALID),
    .m_axi_AWADDR(m_axi_in_13_AWADDR),
    .m_axi_AWBURST(m_axi_in_13_AWBURST),
    .m_axi_AWCACHE(m_axi_in_13_AWCACHE),
    .m_axi_AWID(m_axi_in_13_AWID),
    .m_axi_AWLEN(m_axi_in_13_AWLEN),
    .m_axi_AWLOCK(m_axi_in_13_AWLOCK),
    .m_axi_AWPROT(m_axi_in_13_AWPROT),
    .m_axi_AWQOS(m_axi_in_13_AWQOS),
    .m_axi_AWREADY(m_axi_in_13_AWREADY),
    .m_axi_AWSIZE(m_axi_in_13_AWSIZE),
    .m_axi_AWVALID(m_axi_in_13_AWVALID),
    .m_axi_BID(m_axi_in_13_BID),
    .m_axi_BREADY(m_axi_in_13_BREADY),
    .m_axi_BRESP(m_axi_in_13_BRESP),
    .m_axi_BVALID(m_axi_in_13_BVALID),
    .m_axi_RDATA(m_axi_in_13_RDATA),
    .m_axi_RID(m_axi_in_13_RID),
    .m_axi_RLAST(m_axi_in_13_RLAST),
    .m_axi_RREADY(m_axi_in_13_RREADY),
    .m_axi_RRESP(m_axi_in_13_RRESP),
    .m_axi_RVALID(m_axi_in_13_RVALID),
    .m_axi_WDATA(m_axi_in_13_WDATA),
    .m_axi_WLAST(m_axi_in_13_WLAST),
    .m_axi_WREADY(m_axi_in_13_WREADY),
    .m_axi_WSTRB(m_axi_in_13_WSTRB),
    .m_axi_WVALID(m_axi_in_13_WVALID),
    .read_addr_din(in_13_read_addr__din),
    .read_addr_full_n(in_13_read_addr__full_n),
    .read_addr_write(in_13_read_addr__write),
    .read_data_dout(in_13_read_data__dout),
    .read_data_empty_n(in_13_read_data__empty_n),
    .read_data_read(in_13_read_data__read),
    .write_addr_din(in_13_write_addr__din),
    .write_addr_full_n(in_13_write_addr__full_n),
    .write_addr_write(in_13_write_addr__write),
    .write_data_din(in_13_write_data__din),
    .write_data_full_n(in_13_write_data__full_n),
    .write_data_write(in_13_write_data__write),
    .write_resp_dout(in_13_write_resp__dout),
    .write_resp_empty_n(in_13_write_resp__empty_n),
    .write_resp_read(in_13_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_14__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_14_ARADDR),
    .m_axi_ARBURST(m_axi_in_14_ARBURST),
    .m_axi_ARCACHE(m_axi_in_14_ARCACHE),
    .m_axi_ARID(m_axi_in_14_ARID),
    .m_axi_ARLEN(m_axi_in_14_ARLEN),
    .m_axi_ARLOCK(m_axi_in_14_ARLOCK),
    .m_axi_ARPROT(m_axi_in_14_ARPROT),
    .m_axi_ARQOS(m_axi_in_14_ARQOS),
    .m_axi_ARREADY(m_axi_in_14_ARREADY),
    .m_axi_ARSIZE(m_axi_in_14_ARSIZE),
    .m_axi_ARVALID(m_axi_in_14_ARVALID),
    .m_axi_AWADDR(m_axi_in_14_AWADDR),
    .m_axi_AWBURST(m_axi_in_14_AWBURST),
    .m_axi_AWCACHE(m_axi_in_14_AWCACHE),
    .m_axi_AWID(m_axi_in_14_AWID),
    .m_axi_AWLEN(m_axi_in_14_AWLEN),
    .m_axi_AWLOCK(m_axi_in_14_AWLOCK),
    .m_axi_AWPROT(m_axi_in_14_AWPROT),
    .m_axi_AWQOS(m_axi_in_14_AWQOS),
    .m_axi_AWREADY(m_axi_in_14_AWREADY),
    .m_axi_AWSIZE(m_axi_in_14_AWSIZE),
    .m_axi_AWVALID(m_axi_in_14_AWVALID),
    .m_axi_BID(m_axi_in_14_BID),
    .m_axi_BREADY(m_axi_in_14_BREADY),
    .m_axi_BRESP(m_axi_in_14_BRESP),
    .m_axi_BVALID(m_axi_in_14_BVALID),
    .m_axi_RDATA(m_axi_in_14_RDATA),
    .m_axi_RID(m_axi_in_14_RID),
    .m_axi_RLAST(m_axi_in_14_RLAST),
    .m_axi_RREADY(m_axi_in_14_RREADY),
    .m_axi_RRESP(m_axi_in_14_RRESP),
    .m_axi_RVALID(m_axi_in_14_RVALID),
    .m_axi_WDATA(m_axi_in_14_WDATA),
    .m_axi_WLAST(m_axi_in_14_WLAST),
    .m_axi_WREADY(m_axi_in_14_WREADY),
    .m_axi_WSTRB(m_axi_in_14_WSTRB),
    .m_axi_WVALID(m_axi_in_14_WVALID),
    .read_addr_din(in_14_read_addr__din),
    .read_addr_full_n(in_14_read_addr__full_n),
    .read_addr_write(in_14_read_addr__write),
    .read_data_dout(in_14_read_data__dout),
    .read_data_empty_n(in_14_read_data__empty_n),
    .read_data_read(in_14_read_data__read),
    .write_addr_din(in_14_write_addr__din),
    .write_addr_full_n(in_14_write_addr__full_n),
    .write_addr_write(in_14_write_addr__write),
    .write_data_din(in_14_write_data__din),
    .write_data_full_n(in_14_write_data__full_n),
    .write_data_write(in_14_write_data__write),
    .write_resp_dout(in_14_write_resp__dout),
    .write_resp_empty_n(in_14_write_resp__empty_n),
    .write_resp_read(in_14_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_15__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_15_ARADDR),
    .m_axi_ARBURST(m_axi_in_15_ARBURST),
    .m_axi_ARCACHE(m_axi_in_15_ARCACHE),
    .m_axi_ARID(m_axi_in_15_ARID),
    .m_axi_ARLEN(m_axi_in_15_ARLEN),
    .m_axi_ARLOCK(m_axi_in_15_ARLOCK),
    .m_axi_ARPROT(m_axi_in_15_ARPROT),
    .m_axi_ARQOS(m_axi_in_15_ARQOS),
    .m_axi_ARREADY(m_axi_in_15_ARREADY),
    .m_axi_ARSIZE(m_axi_in_15_ARSIZE),
    .m_axi_ARVALID(m_axi_in_15_ARVALID),
    .m_axi_AWADDR(m_axi_in_15_AWADDR),
    .m_axi_AWBURST(m_axi_in_15_AWBURST),
    .m_axi_AWCACHE(m_axi_in_15_AWCACHE),
    .m_axi_AWID(m_axi_in_15_AWID),
    .m_axi_AWLEN(m_axi_in_15_AWLEN),
    .m_axi_AWLOCK(m_axi_in_15_AWLOCK),
    .m_axi_AWPROT(m_axi_in_15_AWPROT),
    .m_axi_AWQOS(m_axi_in_15_AWQOS),
    .m_axi_AWREADY(m_axi_in_15_AWREADY),
    .m_axi_AWSIZE(m_axi_in_15_AWSIZE),
    .m_axi_AWVALID(m_axi_in_15_AWVALID),
    .m_axi_BID(m_axi_in_15_BID),
    .m_axi_BREADY(m_axi_in_15_BREADY),
    .m_axi_BRESP(m_axi_in_15_BRESP),
    .m_axi_BVALID(m_axi_in_15_BVALID),
    .m_axi_RDATA(m_axi_in_15_RDATA),
    .m_axi_RID(m_axi_in_15_RID),
    .m_axi_RLAST(m_axi_in_15_RLAST),
    .m_axi_RREADY(m_axi_in_15_RREADY),
    .m_axi_RRESP(m_axi_in_15_RRESP),
    .m_axi_RVALID(m_axi_in_15_RVALID),
    .m_axi_WDATA(m_axi_in_15_WDATA),
    .m_axi_WLAST(m_axi_in_15_WLAST),
    .m_axi_WREADY(m_axi_in_15_WREADY),
    .m_axi_WSTRB(m_axi_in_15_WSTRB),
    .m_axi_WVALID(m_axi_in_15_WVALID),
    .read_addr_din(in_15_read_addr__din),
    .read_addr_full_n(in_15_read_addr__full_n),
    .read_addr_write(in_15_read_addr__write),
    .read_data_dout(in_15_read_data__dout),
    .read_data_empty_n(in_15_read_data__empty_n),
    .read_data_read(in_15_read_data__read),
    .write_addr_din(in_15_write_addr__din),
    .write_addr_full_n(in_15_write_addr__full_n),
    .write_addr_write(in_15_write_addr__write),
    .write_data_din(in_15_write_data__din),
    .write_data_full_n(in_15_write_data__full_n),
    .write_data_write(in_15_write_data__write),
    .write_resp_dout(in_15_write_resp__dout),
    .write_resp_empty_n(in_15_write_resp__empty_n),
    .write_resp_read(in_15_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_16__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_16_ARADDR),
    .m_axi_ARBURST(m_axi_in_16_ARBURST),
    .m_axi_ARCACHE(m_axi_in_16_ARCACHE),
    .m_axi_ARID(m_axi_in_16_ARID),
    .m_axi_ARLEN(m_axi_in_16_ARLEN),
    .m_axi_ARLOCK(m_axi_in_16_ARLOCK),
    .m_axi_ARPROT(m_axi_in_16_ARPROT),
    .m_axi_ARQOS(m_axi_in_16_ARQOS),
    .m_axi_ARREADY(m_axi_in_16_ARREADY),
    .m_axi_ARSIZE(m_axi_in_16_ARSIZE),
    .m_axi_ARVALID(m_axi_in_16_ARVALID),
    .m_axi_AWADDR(m_axi_in_16_AWADDR),
    .m_axi_AWBURST(m_axi_in_16_AWBURST),
    .m_axi_AWCACHE(m_axi_in_16_AWCACHE),
    .m_axi_AWID(m_axi_in_16_AWID),
    .m_axi_AWLEN(m_axi_in_16_AWLEN),
    .m_axi_AWLOCK(m_axi_in_16_AWLOCK),
    .m_axi_AWPROT(m_axi_in_16_AWPROT),
    .m_axi_AWQOS(m_axi_in_16_AWQOS),
    .m_axi_AWREADY(m_axi_in_16_AWREADY),
    .m_axi_AWSIZE(m_axi_in_16_AWSIZE),
    .m_axi_AWVALID(m_axi_in_16_AWVALID),
    .m_axi_BID(m_axi_in_16_BID),
    .m_axi_BREADY(m_axi_in_16_BREADY),
    .m_axi_BRESP(m_axi_in_16_BRESP),
    .m_axi_BVALID(m_axi_in_16_BVALID),
    .m_axi_RDATA(m_axi_in_16_RDATA),
    .m_axi_RID(m_axi_in_16_RID),
    .m_axi_RLAST(m_axi_in_16_RLAST),
    .m_axi_RREADY(m_axi_in_16_RREADY),
    .m_axi_RRESP(m_axi_in_16_RRESP),
    .m_axi_RVALID(m_axi_in_16_RVALID),
    .m_axi_WDATA(m_axi_in_16_WDATA),
    .m_axi_WLAST(m_axi_in_16_WLAST),
    .m_axi_WREADY(m_axi_in_16_WREADY),
    .m_axi_WSTRB(m_axi_in_16_WSTRB),
    .m_axi_WVALID(m_axi_in_16_WVALID),
    .read_addr_din(in_16_read_addr__din),
    .read_addr_full_n(in_16_read_addr__full_n),
    .read_addr_write(in_16_read_addr__write),
    .read_data_dout(in_16_read_data__dout),
    .read_data_empty_n(in_16_read_data__empty_n),
    .read_data_read(in_16_read_data__read),
    .write_addr_din(in_16_write_addr__din),
    .write_addr_full_n(in_16_write_addr__full_n),
    .write_addr_write(in_16_write_addr__write),
    .write_data_din(in_16_write_data__din),
    .write_data_full_n(in_16_write_data__full_n),
    .write_data_write(in_16_write_data__write),
    .write_resp_dout(in_16_write_resp__dout),
    .write_resp_empty_n(in_16_write_resp__empty_n),
    .write_resp_read(in_16_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_17__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_17_ARADDR),
    .m_axi_ARBURST(m_axi_in_17_ARBURST),
    .m_axi_ARCACHE(m_axi_in_17_ARCACHE),
    .m_axi_ARID(m_axi_in_17_ARID),
    .m_axi_ARLEN(m_axi_in_17_ARLEN),
    .m_axi_ARLOCK(m_axi_in_17_ARLOCK),
    .m_axi_ARPROT(m_axi_in_17_ARPROT),
    .m_axi_ARQOS(m_axi_in_17_ARQOS),
    .m_axi_ARREADY(m_axi_in_17_ARREADY),
    .m_axi_ARSIZE(m_axi_in_17_ARSIZE),
    .m_axi_ARVALID(m_axi_in_17_ARVALID),
    .m_axi_AWADDR(m_axi_in_17_AWADDR),
    .m_axi_AWBURST(m_axi_in_17_AWBURST),
    .m_axi_AWCACHE(m_axi_in_17_AWCACHE),
    .m_axi_AWID(m_axi_in_17_AWID),
    .m_axi_AWLEN(m_axi_in_17_AWLEN),
    .m_axi_AWLOCK(m_axi_in_17_AWLOCK),
    .m_axi_AWPROT(m_axi_in_17_AWPROT),
    .m_axi_AWQOS(m_axi_in_17_AWQOS),
    .m_axi_AWREADY(m_axi_in_17_AWREADY),
    .m_axi_AWSIZE(m_axi_in_17_AWSIZE),
    .m_axi_AWVALID(m_axi_in_17_AWVALID),
    .m_axi_BID(m_axi_in_17_BID),
    .m_axi_BREADY(m_axi_in_17_BREADY),
    .m_axi_BRESP(m_axi_in_17_BRESP),
    .m_axi_BVALID(m_axi_in_17_BVALID),
    .m_axi_RDATA(m_axi_in_17_RDATA),
    .m_axi_RID(m_axi_in_17_RID),
    .m_axi_RLAST(m_axi_in_17_RLAST),
    .m_axi_RREADY(m_axi_in_17_RREADY),
    .m_axi_RRESP(m_axi_in_17_RRESP),
    .m_axi_RVALID(m_axi_in_17_RVALID),
    .m_axi_WDATA(m_axi_in_17_WDATA),
    .m_axi_WLAST(m_axi_in_17_WLAST),
    .m_axi_WREADY(m_axi_in_17_WREADY),
    .m_axi_WSTRB(m_axi_in_17_WSTRB),
    .m_axi_WVALID(m_axi_in_17_WVALID),
    .read_addr_din(in_17_read_addr__din),
    .read_addr_full_n(in_17_read_addr__full_n),
    .read_addr_write(in_17_read_addr__write),
    .read_data_dout(in_17_read_data__dout),
    .read_data_empty_n(in_17_read_data__empty_n),
    .read_data_read(in_17_read_data__read),
    .write_addr_din(in_17_write_addr__din),
    .write_addr_full_n(in_17_write_addr__full_n),
    .write_addr_write(in_17_write_addr__write),
    .write_data_din(in_17_write_data__din),
    .write_data_full_n(in_17_write_data__full_n),
    .write_data_write(in_17_write_data__write),
    .write_resp_dout(in_17_write_resp__dout),
    .write_resp_empty_n(in_17_write_resp__empty_n),
    .write_resp_read(in_17_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_18__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_18_ARADDR),
    .m_axi_ARBURST(m_axi_in_18_ARBURST),
    .m_axi_ARCACHE(m_axi_in_18_ARCACHE),
    .m_axi_ARID(m_axi_in_18_ARID),
    .m_axi_ARLEN(m_axi_in_18_ARLEN),
    .m_axi_ARLOCK(m_axi_in_18_ARLOCK),
    .m_axi_ARPROT(m_axi_in_18_ARPROT),
    .m_axi_ARQOS(m_axi_in_18_ARQOS),
    .m_axi_ARREADY(m_axi_in_18_ARREADY),
    .m_axi_ARSIZE(m_axi_in_18_ARSIZE),
    .m_axi_ARVALID(m_axi_in_18_ARVALID),
    .m_axi_AWADDR(m_axi_in_18_AWADDR),
    .m_axi_AWBURST(m_axi_in_18_AWBURST),
    .m_axi_AWCACHE(m_axi_in_18_AWCACHE),
    .m_axi_AWID(m_axi_in_18_AWID),
    .m_axi_AWLEN(m_axi_in_18_AWLEN),
    .m_axi_AWLOCK(m_axi_in_18_AWLOCK),
    .m_axi_AWPROT(m_axi_in_18_AWPROT),
    .m_axi_AWQOS(m_axi_in_18_AWQOS),
    .m_axi_AWREADY(m_axi_in_18_AWREADY),
    .m_axi_AWSIZE(m_axi_in_18_AWSIZE),
    .m_axi_AWVALID(m_axi_in_18_AWVALID),
    .m_axi_BID(m_axi_in_18_BID),
    .m_axi_BREADY(m_axi_in_18_BREADY),
    .m_axi_BRESP(m_axi_in_18_BRESP),
    .m_axi_BVALID(m_axi_in_18_BVALID),
    .m_axi_RDATA(m_axi_in_18_RDATA),
    .m_axi_RID(m_axi_in_18_RID),
    .m_axi_RLAST(m_axi_in_18_RLAST),
    .m_axi_RREADY(m_axi_in_18_RREADY),
    .m_axi_RRESP(m_axi_in_18_RRESP),
    .m_axi_RVALID(m_axi_in_18_RVALID),
    .m_axi_WDATA(m_axi_in_18_WDATA),
    .m_axi_WLAST(m_axi_in_18_WLAST),
    .m_axi_WREADY(m_axi_in_18_WREADY),
    .m_axi_WSTRB(m_axi_in_18_WSTRB),
    .m_axi_WVALID(m_axi_in_18_WVALID),
    .read_addr_din(in_18_read_addr__din),
    .read_addr_full_n(in_18_read_addr__full_n),
    .read_addr_write(in_18_read_addr__write),
    .read_data_dout(in_18_read_data__dout),
    .read_data_empty_n(in_18_read_data__empty_n),
    .read_data_read(in_18_read_data__read),
    .write_addr_din(in_18_write_addr__din),
    .write_addr_full_n(in_18_write_addr__full_n),
    .write_addr_write(in_18_write_addr__write),
    .write_data_din(in_18_write_data__din),
    .write_data_full_n(in_18_write_data__full_n),
    .write_data_write(in_18_write_data__write),
    .write_resp_dout(in_18_write_resp__dout),
    .write_resp_empty_n(in_18_write_resp__empty_n),
    .write_resp_read(in_18_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_19__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_19_ARADDR),
    .m_axi_ARBURST(m_axi_in_19_ARBURST),
    .m_axi_ARCACHE(m_axi_in_19_ARCACHE),
    .m_axi_ARID(m_axi_in_19_ARID),
    .m_axi_ARLEN(m_axi_in_19_ARLEN),
    .m_axi_ARLOCK(m_axi_in_19_ARLOCK),
    .m_axi_ARPROT(m_axi_in_19_ARPROT),
    .m_axi_ARQOS(m_axi_in_19_ARQOS),
    .m_axi_ARREADY(m_axi_in_19_ARREADY),
    .m_axi_ARSIZE(m_axi_in_19_ARSIZE),
    .m_axi_ARVALID(m_axi_in_19_ARVALID),
    .m_axi_AWADDR(m_axi_in_19_AWADDR),
    .m_axi_AWBURST(m_axi_in_19_AWBURST),
    .m_axi_AWCACHE(m_axi_in_19_AWCACHE),
    .m_axi_AWID(m_axi_in_19_AWID),
    .m_axi_AWLEN(m_axi_in_19_AWLEN),
    .m_axi_AWLOCK(m_axi_in_19_AWLOCK),
    .m_axi_AWPROT(m_axi_in_19_AWPROT),
    .m_axi_AWQOS(m_axi_in_19_AWQOS),
    .m_axi_AWREADY(m_axi_in_19_AWREADY),
    .m_axi_AWSIZE(m_axi_in_19_AWSIZE),
    .m_axi_AWVALID(m_axi_in_19_AWVALID),
    .m_axi_BID(m_axi_in_19_BID),
    .m_axi_BREADY(m_axi_in_19_BREADY),
    .m_axi_BRESP(m_axi_in_19_BRESP),
    .m_axi_BVALID(m_axi_in_19_BVALID),
    .m_axi_RDATA(m_axi_in_19_RDATA),
    .m_axi_RID(m_axi_in_19_RID),
    .m_axi_RLAST(m_axi_in_19_RLAST),
    .m_axi_RREADY(m_axi_in_19_RREADY),
    .m_axi_RRESP(m_axi_in_19_RRESP),
    .m_axi_RVALID(m_axi_in_19_RVALID),
    .m_axi_WDATA(m_axi_in_19_WDATA),
    .m_axi_WLAST(m_axi_in_19_WLAST),
    .m_axi_WREADY(m_axi_in_19_WREADY),
    .m_axi_WSTRB(m_axi_in_19_WSTRB),
    .m_axi_WVALID(m_axi_in_19_WVALID),
    .read_addr_din(in_19_read_addr__din),
    .read_addr_full_n(in_19_read_addr__full_n),
    .read_addr_write(in_19_read_addr__write),
    .read_data_dout(in_19_read_data__dout),
    .read_data_empty_n(in_19_read_data__empty_n),
    .read_data_read(in_19_read_data__read),
    .write_addr_din(in_19_write_addr__din),
    .write_addr_full_n(in_19_write_addr__full_n),
    .write_addr_write(in_19_write_addr__write),
    .write_data_din(in_19_write_data__din),
    .write_data_full_n(in_19_write_data__full_n),
    .write_data_write(in_19_write_data__write),
    .write_resp_dout(in_19_write_resp__dout),
    .write_resp_empty_n(in_19_write_resp__empty_n),
    .write_resp_read(in_19_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_2_ARADDR),
    .m_axi_ARBURST(m_axi_in_2_ARBURST),
    .m_axi_ARCACHE(m_axi_in_2_ARCACHE),
    .m_axi_ARID(m_axi_in_2_ARID),
    .m_axi_ARLEN(m_axi_in_2_ARLEN),
    .m_axi_ARLOCK(m_axi_in_2_ARLOCK),
    .m_axi_ARPROT(m_axi_in_2_ARPROT),
    .m_axi_ARQOS(m_axi_in_2_ARQOS),
    .m_axi_ARREADY(m_axi_in_2_ARREADY),
    .m_axi_ARSIZE(m_axi_in_2_ARSIZE),
    .m_axi_ARVALID(m_axi_in_2_ARVALID),
    .m_axi_AWADDR(m_axi_in_2_AWADDR),
    .m_axi_AWBURST(m_axi_in_2_AWBURST),
    .m_axi_AWCACHE(m_axi_in_2_AWCACHE),
    .m_axi_AWID(m_axi_in_2_AWID),
    .m_axi_AWLEN(m_axi_in_2_AWLEN),
    .m_axi_AWLOCK(m_axi_in_2_AWLOCK),
    .m_axi_AWPROT(m_axi_in_2_AWPROT),
    .m_axi_AWQOS(m_axi_in_2_AWQOS),
    .m_axi_AWREADY(m_axi_in_2_AWREADY),
    .m_axi_AWSIZE(m_axi_in_2_AWSIZE),
    .m_axi_AWVALID(m_axi_in_2_AWVALID),
    .m_axi_BID(m_axi_in_2_BID),
    .m_axi_BREADY(m_axi_in_2_BREADY),
    .m_axi_BRESP(m_axi_in_2_BRESP),
    .m_axi_BVALID(m_axi_in_2_BVALID),
    .m_axi_RDATA(m_axi_in_2_RDATA),
    .m_axi_RID(m_axi_in_2_RID),
    .m_axi_RLAST(m_axi_in_2_RLAST),
    .m_axi_RREADY(m_axi_in_2_RREADY),
    .m_axi_RRESP(m_axi_in_2_RRESP),
    .m_axi_RVALID(m_axi_in_2_RVALID),
    .m_axi_WDATA(m_axi_in_2_WDATA),
    .m_axi_WLAST(m_axi_in_2_WLAST),
    .m_axi_WREADY(m_axi_in_2_WREADY),
    .m_axi_WSTRB(m_axi_in_2_WSTRB),
    .m_axi_WVALID(m_axi_in_2_WVALID),
    .read_addr_din(in_2_read_addr__din),
    .read_addr_full_n(in_2_read_addr__full_n),
    .read_addr_write(in_2_read_addr__write),
    .read_data_dout(in_2_read_data__dout),
    .read_data_empty_n(in_2_read_data__empty_n),
    .read_data_read(in_2_read_data__read),
    .write_addr_din(in_2_write_addr__din),
    .write_addr_full_n(in_2_write_addr__full_n),
    .write_addr_write(in_2_write_addr__write),
    .write_data_din(in_2_write_data__din),
    .write_data_full_n(in_2_write_data__full_n),
    .write_data_write(in_2_write_data__write),
    .write_resp_dout(in_2_write_resp__dout),
    .write_resp_empty_n(in_2_write_resp__empty_n),
    .write_resp_read(in_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_20__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_20_ARADDR),
    .m_axi_ARBURST(m_axi_in_20_ARBURST),
    .m_axi_ARCACHE(m_axi_in_20_ARCACHE),
    .m_axi_ARID(m_axi_in_20_ARID),
    .m_axi_ARLEN(m_axi_in_20_ARLEN),
    .m_axi_ARLOCK(m_axi_in_20_ARLOCK),
    .m_axi_ARPROT(m_axi_in_20_ARPROT),
    .m_axi_ARQOS(m_axi_in_20_ARQOS),
    .m_axi_ARREADY(m_axi_in_20_ARREADY),
    .m_axi_ARSIZE(m_axi_in_20_ARSIZE),
    .m_axi_ARVALID(m_axi_in_20_ARVALID),
    .m_axi_AWADDR(m_axi_in_20_AWADDR),
    .m_axi_AWBURST(m_axi_in_20_AWBURST),
    .m_axi_AWCACHE(m_axi_in_20_AWCACHE),
    .m_axi_AWID(m_axi_in_20_AWID),
    .m_axi_AWLEN(m_axi_in_20_AWLEN),
    .m_axi_AWLOCK(m_axi_in_20_AWLOCK),
    .m_axi_AWPROT(m_axi_in_20_AWPROT),
    .m_axi_AWQOS(m_axi_in_20_AWQOS),
    .m_axi_AWREADY(m_axi_in_20_AWREADY),
    .m_axi_AWSIZE(m_axi_in_20_AWSIZE),
    .m_axi_AWVALID(m_axi_in_20_AWVALID),
    .m_axi_BID(m_axi_in_20_BID),
    .m_axi_BREADY(m_axi_in_20_BREADY),
    .m_axi_BRESP(m_axi_in_20_BRESP),
    .m_axi_BVALID(m_axi_in_20_BVALID),
    .m_axi_RDATA(m_axi_in_20_RDATA),
    .m_axi_RID(m_axi_in_20_RID),
    .m_axi_RLAST(m_axi_in_20_RLAST),
    .m_axi_RREADY(m_axi_in_20_RREADY),
    .m_axi_RRESP(m_axi_in_20_RRESP),
    .m_axi_RVALID(m_axi_in_20_RVALID),
    .m_axi_WDATA(m_axi_in_20_WDATA),
    .m_axi_WLAST(m_axi_in_20_WLAST),
    .m_axi_WREADY(m_axi_in_20_WREADY),
    .m_axi_WSTRB(m_axi_in_20_WSTRB),
    .m_axi_WVALID(m_axi_in_20_WVALID),
    .read_addr_din(in_20_read_addr__din),
    .read_addr_full_n(in_20_read_addr__full_n),
    .read_addr_write(in_20_read_addr__write),
    .read_data_dout(in_20_read_data__dout),
    .read_data_empty_n(in_20_read_data__empty_n),
    .read_data_read(in_20_read_data__read),
    .write_addr_din(in_20_write_addr__din),
    .write_addr_full_n(in_20_write_addr__full_n),
    .write_addr_write(in_20_write_addr__write),
    .write_data_din(in_20_write_data__din),
    .write_data_full_n(in_20_write_data__full_n),
    .write_data_write(in_20_write_data__write),
    .write_resp_dout(in_20_write_resp__dout),
    .write_resp_empty_n(in_20_write_resp__empty_n),
    .write_resp_read(in_20_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_21__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_21_ARADDR),
    .m_axi_ARBURST(m_axi_in_21_ARBURST),
    .m_axi_ARCACHE(m_axi_in_21_ARCACHE),
    .m_axi_ARID(m_axi_in_21_ARID),
    .m_axi_ARLEN(m_axi_in_21_ARLEN),
    .m_axi_ARLOCK(m_axi_in_21_ARLOCK),
    .m_axi_ARPROT(m_axi_in_21_ARPROT),
    .m_axi_ARQOS(m_axi_in_21_ARQOS),
    .m_axi_ARREADY(m_axi_in_21_ARREADY),
    .m_axi_ARSIZE(m_axi_in_21_ARSIZE),
    .m_axi_ARVALID(m_axi_in_21_ARVALID),
    .m_axi_AWADDR(m_axi_in_21_AWADDR),
    .m_axi_AWBURST(m_axi_in_21_AWBURST),
    .m_axi_AWCACHE(m_axi_in_21_AWCACHE),
    .m_axi_AWID(m_axi_in_21_AWID),
    .m_axi_AWLEN(m_axi_in_21_AWLEN),
    .m_axi_AWLOCK(m_axi_in_21_AWLOCK),
    .m_axi_AWPROT(m_axi_in_21_AWPROT),
    .m_axi_AWQOS(m_axi_in_21_AWQOS),
    .m_axi_AWREADY(m_axi_in_21_AWREADY),
    .m_axi_AWSIZE(m_axi_in_21_AWSIZE),
    .m_axi_AWVALID(m_axi_in_21_AWVALID),
    .m_axi_BID(m_axi_in_21_BID),
    .m_axi_BREADY(m_axi_in_21_BREADY),
    .m_axi_BRESP(m_axi_in_21_BRESP),
    .m_axi_BVALID(m_axi_in_21_BVALID),
    .m_axi_RDATA(m_axi_in_21_RDATA),
    .m_axi_RID(m_axi_in_21_RID),
    .m_axi_RLAST(m_axi_in_21_RLAST),
    .m_axi_RREADY(m_axi_in_21_RREADY),
    .m_axi_RRESP(m_axi_in_21_RRESP),
    .m_axi_RVALID(m_axi_in_21_RVALID),
    .m_axi_WDATA(m_axi_in_21_WDATA),
    .m_axi_WLAST(m_axi_in_21_WLAST),
    .m_axi_WREADY(m_axi_in_21_WREADY),
    .m_axi_WSTRB(m_axi_in_21_WSTRB),
    .m_axi_WVALID(m_axi_in_21_WVALID),
    .read_addr_din(in_21_read_addr__din),
    .read_addr_full_n(in_21_read_addr__full_n),
    .read_addr_write(in_21_read_addr__write),
    .read_data_dout(in_21_read_data__dout),
    .read_data_empty_n(in_21_read_data__empty_n),
    .read_data_read(in_21_read_data__read),
    .write_addr_din(in_21_write_addr__din),
    .write_addr_full_n(in_21_write_addr__full_n),
    .write_addr_write(in_21_write_addr__write),
    .write_data_din(in_21_write_data__din),
    .write_data_full_n(in_21_write_data__full_n),
    .write_data_write(in_21_write_data__write),
    .write_resp_dout(in_21_write_resp__dout),
    .write_resp_empty_n(in_21_write_resp__empty_n),
    .write_resp_read(in_21_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_22__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_22_ARADDR),
    .m_axi_ARBURST(m_axi_in_22_ARBURST),
    .m_axi_ARCACHE(m_axi_in_22_ARCACHE),
    .m_axi_ARID(m_axi_in_22_ARID),
    .m_axi_ARLEN(m_axi_in_22_ARLEN),
    .m_axi_ARLOCK(m_axi_in_22_ARLOCK),
    .m_axi_ARPROT(m_axi_in_22_ARPROT),
    .m_axi_ARQOS(m_axi_in_22_ARQOS),
    .m_axi_ARREADY(m_axi_in_22_ARREADY),
    .m_axi_ARSIZE(m_axi_in_22_ARSIZE),
    .m_axi_ARVALID(m_axi_in_22_ARVALID),
    .m_axi_AWADDR(m_axi_in_22_AWADDR),
    .m_axi_AWBURST(m_axi_in_22_AWBURST),
    .m_axi_AWCACHE(m_axi_in_22_AWCACHE),
    .m_axi_AWID(m_axi_in_22_AWID),
    .m_axi_AWLEN(m_axi_in_22_AWLEN),
    .m_axi_AWLOCK(m_axi_in_22_AWLOCK),
    .m_axi_AWPROT(m_axi_in_22_AWPROT),
    .m_axi_AWQOS(m_axi_in_22_AWQOS),
    .m_axi_AWREADY(m_axi_in_22_AWREADY),
    .m_axi_AWSIZE(m_axi_in_22_AWSIZE),
    .m_axi_AWVALID(m_axi_in_22_AWVALID),
    .m_axi_BID(m_axi_in_22_BID),
    .m_axi_BREADY(m_axi_in_22_BREADY),
    .m_axi_BRESP(m_axi_in_22_BRESP),
    .m_axi_BVALID(m_axi_in_22_BVALID),
    .m_axi_RDATA(m_axi_in_22_RDATA),
    .m_axi_RID(m_axi_in_22_RID),
    .m_axi_RLAST(m_axi_in_22_RLAST),
    .m_axi_RREADY(m_axi_in_22_RREADY),
    .m_axi_RRESP(m_axi_in_22_RRESP),
    .m_axi_RVALID(m_axi_in_22_RVALID),
    .m_axi_WDATA(m_axi_in_22_WDATA),
    .m_axi_WLAST(m_axi_in_22_WLAST),
    .m_axi_WREADY(m_axi_in_22_WREADY),
    .m_axi_WSTRB(m_axi_in_22_WSTRB),
    .m_axi_WVALID(m_axi_in_22_WVALID),
    .read_addr_din(in_22_read_addr__din),
    .read_addr_full_n(in_22_read_addr__full_n),
    .read_addr_write(in_22_read_addr__write),
    .read_data_dout(in_22_read_data__dout),
    .read_data_empty_n(in_22_read_data__empty_n),
    .read_data_read(in_22_read_data__read),
    .write_addr_din(in_22_write_addr__din),
    .write_addr_full_n(in_22_write_addr__full_n),
    .write_addr_write(in_22_write_addr__write),
    .write_data_din(in_22_write_data__din),
    .write_data_full_n(in_22_write_data__full_n),
    .write_data_write(in_22_write_data__write),
    .write_resp_dout(in_22_write_resp__dout),
    .write_resp_empty_n(in_22_write_resp__empty_n),
    .write_resp_read(in_22_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_23__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_23_ARADDR),
    .m_axi_ARBURST(m_axi_in_23_ARBURST),
    .m_axi_ARCACHE(m_axi_in_23_ARCACHE),
    .m_axi_ARID(m_axi_in_23_ARID),
    .m_axi_ARLEN(m_axi_in_23_ARLEN),
    .m_axi_ARLOCK(m_axi_in_23_ARLOCK),
    .m_axi_ARPROT(m_axi_in_23_ARPROT),
    .m_axi_ARQOS(m_axi_in_23_ARQOS),
    .m_axi_ARREADY(m_axi_in_23_ARREADY),
    .m_axi_ARSIZE(m_axi_in_23_ARSIZE),
    .m_axi_ARVALID(m_axi_in_23_ARVALID),
    .m_axi_AWADDR(m_axi_in_23_AWADDR),
    .m_axi_AWBURST(m_axi_in_23_AWBURST),
    .m_axi_AWCACHE(m_axi_in_23_AWCACHE),
    .m_axi_AWID(m_axi_in_23_AWID),
    .m_axi_AWLEN(m_axi_in_23_AWLEN),
    .m_axi_AWLOCK(m_axi_in_23_AWLOCK),
    .m_axi_AWPROT(m_axi_in_23_AWPROT),
    .m_axi_AWQOS(m_axi_in_23_AWQOS),
    .m_axi_AWREADY(m_axi_in_23_AWREADY),
    .m_axi_AWSIZE(m_axi_in_23_AWSIZE),
    .m_axi_AWVALID(m_axi_in_23_AWVALID),
    .m_axi_BID(m_axi_in_23_BID),
    .m_axi_BREADY(m_axi_in_23_BREADY),
    .m_axi_BRESP(m_axi_in_23_BRESP),
    .m_axi_BVALID(m_axi_in_23_BVALID),
    .m_axi_RDATA(m_axi_in_23_RDATA),
    .m_axi_RID(m_axi_in_23_RID),
    .m_axi_RLAST(m_axi_in_23_RLAST),
    .m_axi_RREADY(m_axi_in_23_RREADY),
    .m_axi_RRESP(m_axi_in_23_RRESP),
    .m_axi_RVALID(m_axi_in_23_RVALID),
    .m_axi_WDATA(m_axi_in_23_WDATA),
    .m_axi_WLAST(m_axi_in_23_WLAST),
    .m_axi_WREADY(m_axi_in_23_WREADY),
    .m_axi_WSTRB(m_axi_in_23_WSTRB),
    .m_axi_WVALID(m_axi_in_23_WVALID),
    .read_addr_din(in_23_read_addr__din),
    .read_addr_full_n(in_23_read_addr__full_n),
    .read_addr_write(in_23_read_addr__write),
    .read_data_dout(in_23_read_data__dout),
    .read_data_empty_n(in_23_read_data__empty_n),
    .read_data_read(in_23_read_data__read),
    .write_addr_din(in_23_write_addr__din),
    .write_addr_full_n(in_23_write_addr__full_n),
    .write_addr_write(in_23_write_addr__write),
    .write_data_din(in_23_write_data__din),
    .write_data_full_n(in_23_write_data__full_n),
    .write_data_write(in_23_write_data__write),
    .write_resp_dout(in_23_write_resp__dout),
    .write_resp_empty_n(in_23_write_resp__empty_n),
    .write_resp_read(in_23_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_24__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_24_ARADDR),
    .m_axi_ARBURST(m_axi_in_24_ARBURST),
    .m_axi_ARCACHE(m_axi_in_24_ARCACHE),
    .m_axi_ARID(m_axi_in_24_ARID),
    .m_axi_ARLEN(m_axi_in_24_ARLEN),
    .m_axi_ARLOCK(m_axi_in_24_ARLOCK),
    .m_axi_ARPROT(m_axi_in_24_ARPROT),
    .m_axi_ARQOS(m_axi_in_24_ARQOS),
    .m_axi_ARREADY(m_axi_in_24_ARREADY),
    .m_axi_ARSIZE(m_axi_in_24_ARSIZE),
    .m_axi_ARVALID(m_axi_in_24_ARVALID),
    .m_axi_AWADDR(m_axi_in_24_AWADDR),
    .m_axi_AWBURST(m_axi_in_24_AWBURST),
    .m_axi_AWCACHE(m_axi_in_24_AWCACHE),
    .m_axi_AWID(m_axi_in_24_AWID),
    .m_axi_AWLEN(m_axi_in_24_AWLEN),
    .m_axi_AWLOCK(m_axi_in_24_AWLOCK),
    .m_axi_AWPROT(m_axi_in_24_AWPROT),
    .m_axi_AWQOS(m_axi_in_24_AWQOS),
    .m_axi_AWREADY(m_axi_in_24_AWREADY),
    .m_axi_AWSIZE(m_axi_in_24_AWSIZE),
    .m_axi_AWVALID(m_axi_in_24_AWVALID),
    .m_axi_BID(m_axi_in_24_BID),
    .m_axi_BREADY(m_axi_in_24_BREADY),
    .m_axi_BRESP(m_axi_in_24_BRESP),
    .m_axi_BVALID(m_axi_in_24_BVALID),
    .m_axi_RDATA(m_axi_in_24_RDATA),
    .m_axi_RID(m_axi_in_24_RID),
    .m_axi_RLAST(m_axi_in_24_RLAST),
    .m_axi_RREADY(m_axi_in_24_RREADY),
    .m_axi_RRESP(m_axi_in_24_RRESP),
    .m_axi_RVALID(m_axi_in_24_RVALID),
    .m_axi_WDATA(m_axi_in_24_WDATA),
    .m_axi_WLAST(m_axi_in_24_WLAST),
    .m_axi_WREADY(m_axi_in_24_WREADY),
    .m_axi_WSTRB(m_axi_in_24_WSTRB),
    .m_axi_WVALID(m_axi_in_24_WVALID),
    .read_addr_din(in_24_read_addr__din),
    .read_addr_full_n(in_24_read_addr__full_n),
    .read_addr_write(in_24_read_addr__write),
    .read_data_dout(in_24_read_data__dout),
    .read_data_empty_n(in_24_read_data__empty_n),
    .read_data_read(in_24_read_data__read),
    .write_addr_din(in_24_write_addr__din),
    .write_addr_full_n(in_24_write_addr__full_n),
    .write_addr_write(in_24_write_addr__write),
    .write_data_din(in_24_write_data__din),
    .write_data_full_n(in_24_write_data__full_n),
    .write_data_write(in_24_write_data__write),
    .write_resp_dout(in_24_write_resp__dout),
    .write_resp_empty_n(in_24_write_resp__empty_n),
    .write_resp_read(in_24_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_25__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_25_ARADDR),
    .m_axi_ARBURST(m_axi_in_25_ARBURST),
    .m_axi_ARCACHE(m_axi_in_25_ARCACHE),
    .m_axi_ARID(m_axi_in_25_ARID),
    .m_axi_ARLEN(m_axi_in_25_ARLEN),
    .m_axi_ARLOCK(m_axi_in_25_ARLOCK),
    .m_axi_ARPROT(m_axi_in_25_ARPROT),
    .m_axi_ARQOS(m_axi_in_25_ARQOS),
    .m_axi_ARREADY(m_axi_in_25_ARREADY),
    .m_axi_ARSIZE(m_axi_in_25_ARSIZE),
    .m_axi_ARVALID(m_axi_in_25_ARVALID),
    .m_axi_AWADDR(m_axi_in_25_AWADDR),
    .m_axi_AWBURST(m_axi_in_25_AWBURST),
    .m_axi_AWCACHE(m_axi_in_25_AWCACHE),
    .m_axi_AWID(m_axi_in_25_AWID),
    .m_axi_AWLEN(m_axi_in_25_AWLEN),
    .m_axi_AWLOCK(m_axi_in_25_AWLOCK),
    .m_axi_AWPROT(m_axi_in_25_AWPROT),
    .m_axi_AWQOS(m_axi_in_25_AWQOS),
    .m_axi_AWREADY(m_axi_in_25_AWREADY),
    .m_axi_AWSIZE(m_axi_in_25_AWSIZE),
    .m_axi_AWVALID(m_axi_in_25_AWVALID),
    .m_axi_BID(m_axi_in_25_BID),
    .m_axi_BREADY(m_axi_in_25_BREADY),
    .m_axi_BRESP(m_axi_in_25_BRESP),
    .m_axi_BVALID(m_axi_in_25_BVALID),
    .m_axi_RDATA(m_axi_in_25_RDATA),
    .m_axi_RID(m_axi_in_25_RID),
    .m_axi_RLAST(m_axi_in_25_RLAST),
    .m_axi_RREADY(m_axi_in_25_RREADY),
    .m_axi_RRESP(m_axi_in_25_RRESP),
    .m_axi_RVALID(m_axi_in_25_RVALID),
    .m_axi_WDATA(m_axi_in_25_WDATA),
    .m_axi_WLAST(m_axi_in_25_WLAST),
    .m_axi_WREADY(m_axi_in_25_WREADY),
    .m_axi_WSTRB(m_axi_in_25_WSTRB),
    .m_axi_WVALID(m_axi_in_25_WVALID),
    .read_addr_din(in_25_read_addr__din),
    .read_addr_full_n(in_25_read_addr__full_n),
    .read_addr_write(in_25_read_addr__write),
    .read_data_dout(in_25_read_data__dout),
    .read_data_empty_n(in_25_read_data__empty_n),
    .read_data_read(in_25_read_data__read),
    .write_addr_din(in_25_write_addr__din),
    .write_addr_full_n(in_25_write_addr__full_n),
    .write_addr_write(in_25_write_addr__write),
    .write_data_din(in_25_write_data__din),
    .write_data_full_n(in_25_write_data__full_n),
    .write_data_write(in_25_write_data__write),
    .write_resp_dout(in_25_write_resp__dout),
    .write_resp_empty_n(in_25_write_resp__empty_n),
    .write_resp_read(in_25_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_26__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_26_ARADDR),
    .m_axi_ARBURST(m_axi_in_26_ARBURST),
    .m_axi_ARCACHE(m_axi_in_26_ARCACHE),
    .m_axi_ARID(m_axi_in_26_ARID),
    .m_axi_ARLEN(m_axi_in_26_ARLEN),
    .m_axi_ARLOCK(m_axi_in_26_ARLOCK),
    .m_axi_ARPROT(m_axi_in_26_ARPROT),
    .m_axi_ARQOS(m_axi_in_26_ARQOS),
    .m_axi_ARREADY(m_axi_in_26_ARREADY),
    .m_axi_ARSIZE(m_axi_in_26_ARSIZE),
    .m_axi_ARVALID(m_axi_in_26_ARVALID),
    .m_axi_AWADDR(m_axi_in_26_AWADDR),
    .m_axi_AWBURST(m_axi_in_26_AWBURST),
    .m_axi_AWCACHE(m_axi_in_26_AWCACHE),
    .m_axi_AWID(m_axi_in_26_AWID),
    .m_axi_AWLEN(m_axi_in_26_AWLEN),
    .m_axi_AWLOCK(m_axi_in_26_AWLOCK),
    .m_axi_AWPROT(m_axi_in_26_AWPROT),
    .m_axi_AWQOS(m_axi_in_26_AWQOS),
    .m_axi_AWREADY(m_axi_in_26_AWREADY),
    .m_axi_AWSIZE(m_axi_in_26_AWSIZE),
    .m_axi_AWVALID(m_axi_in_26_AWVALID),
    .m_axi_BID(m_axi_in_26_BID),
    .m_axi_BREADY(m_axi_in_26_BREADY),
    .m_axi_BRESP(m_axi_in_26_BRESP),
    .m_axi_BVALID(m_axi_in_26_BVALID),
    .m_axi_RDATA(m_axi_in_26_RDATA),
    .m_axi_RID(m_axi_in_26_RID),
    .m_axi_RLAST(m_axi_in_26_RLAST),
    .m_axi_RREADY(m_axi_in_26_RREADY),
    .m_axi_RRESP(m_axi_in_26_RRESP),
    .m_axi_RVALID(m_axi_in_26_RVALID),
    .m_axi_WDATA(m_axi_in_26_WDATA),
    .m_axi_WLAST(m_axi_in_26_WLAST),
    .m_axi_WREADY(m_axi_in_26_WREADY),
    .m_axi_WSTRB(m_axi_in_26_WSTRB),
    .m_axi_WVALID(m_axi_in_26_WVALID),
    .read_addr_din(in_26_read_addr__din),
    .read_addr_full_n(in_26_read_addr__full_n),
    .read_addr_write(in_26_read_addr__write),
    .read_data_dout(in_26_read_data__dout),
    .read_data_empty_n(in_26_read_data__empty_n),
    .read_data_read(in_26_read_data__read),
    .write_addr_din(in_26_write_addr__din),
    .write_addr_full_n(in_26_write_addr__full_n),
    .write_addr_write(in_26_write_addr__write),
    .write_data_din(in_26_write_data__din),
    .write_data_full_n(in_26_write_data__full_n),
    .write_data_write(in_26_write_data__write),
    .write_resp_dout(in_26_write_resp__dout),
    .write_resp_empty_n(in_26_write_resp__empty_n),
    .write_resp_read(in_26_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_27__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_27_ARADDR),
    .m_axi_ARBURST(m_axi_in_27_ARBURST),
    .m_axi_ARCACHE(m_axi_in_27_ARCACHE),
    .m_axi_ARID(m_axi_in_27_ARID),
    .m_axi_ARLEN(m_axi_in_27_ARLEN),
    .m_axi_ARLOCK(m_axi_in_27_ARLOCK),
    .m_axi_ARPROT(m_axi_in_27_ARPROT),
    .m_axi_ARQOS(m_axi_in_27_ARQOS),
    .m_axi_ARREADY(m_axi_in_27_ARREADY),
    .m_axi_ARSIZE(m_axi_in_27_ARSIZE),
    .m_axi_ARVALID(m_axi_in_27_ARVALID),
    .m_axi_AWADDR(m_axi_in_27_AWADDR),
    .m_axi_AWBURST(m_axi_in_27_AWBURST),
    .m_axi_AWCACHE(m_axi_in_27_AWCACHE),
    .m_axi_AWID(m_axi_in_27_AWID),
    .m_axi_AWLEN(m_axi_in_27_AWLEN),
    .m_axi_AWLOCK(m_axi_in_27_AWLOCK),
    .m_axi_AWPROT(m_axi_in_27_AWPROT),
    .m_axi_AWQOS(m_axi_in_27_AWQOS),
    .m_axi_AWREADY(m_axi_in_27_AWREADY),
    .m_axi_AWSIZE(m_axi_in_27_AWSIZE),
    .m_axi_AWVALID(m_axi_in_27_AWVALID),
    .m_axi_BID(m_axi_in_27_BID),
    .m_axi_BREADY(m_axi_in_27_BREADY),
    .m_axi_BRESP(m_axi_in_27_BRESP),
    .m_axi_BVALID(m_axi_in_27_BVALID),
    .m_axi_RDATA(m_axi_in_27_RDATA),
    .m_axi_RID(m_axi_in_27_RID),
    .m_axi_RLAST(m_axi_in_27_RLAST),
    .m_axi_RREADY(m_axi_in_27_RREADY),
    .m_axi_RRESP(m_axi_in_27_RRESP),
    .m_axi_RVALID(m_axi_in_27_RVALID),
    .m_axi_WDATA(m_axi_in_27_WDATA),
    .m_axi_WLAST(m_axi_in_27_WLAST),
    .m_axi_WREADY(m_axi_in_27_WREADY),
    .m_axi_WSTRB(m_axi_in_27_WSTRB),
    .m_axi_WVALID(m_axi_in_27_WVALID),
    .read_addr_din(in_27_read_addr__din),
    .read_addr_full_n(in_27_read_addr__full_n),
    .read_addr_write(in_27_read_addr__write),
    .read_data_dout(in_27_read_data__dout),
    .read_data_empty_n(in_27_read_data__empty_n),
    .read_data_read(in_27_read_data__read),
    .write_addr_din(in_27_write_addr__din),
    .write_addr_full_n(in_27_write_addr__full_n),
    .write_addr_write(in_27_write_addr__write),
    .write_data_din(in_27_write_data__din),
    .write_data_full_n(in_27_write_data__full_n),
    .write_data_write(in_27_write_data__write),
    .write_resp_dout(in_27_write_resp__dout),
    .write_resp_empty_n(in_27_write_resp__empty_n),
    .write_resp_read(in_27_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_28__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_28_ARADDR),
    .m_axi_ARBURST(m_axi_in_28_ARBURST),
    .m_axi_ARCACHE(m_axi_in_28_ARCACHE),
    .m_axi_ARID(m_axi_in_28_ARID),
    .m_axi_ARLEN(m_axi_in_28_ARLEN),
    .m_axi_ARLOCK(m_axi_in_28_ARLOCK),
    .m_axi_ARPROT(m_axi_in_28_ARPROT),
    .m_axi_ARQOS(m_axi_in_28_ARQOS),
    .m_axi_ARREADY(m_axi_in_28_ARREADY),
    .m_axi_ARSIZE(m_axi_in_28_ARSIZE),
    .m_axi_ARVALID(m_axi_in_28_ARVALID),
    .m_axi_AWADDR(m_axi_in_28_AWADDR),
    .m_axi_AWBURST(m_axi_in_28_AWBURST),
    .m_axi_AWCACHE(m_axi_in_28_AWCACHE),
    .m_axi_AWID(m_axi_in_28_AWID),
    .m_axi_AWLEN(m_axi_in_28_AWLEN),
    .m_axi_AWLOCK(m_axi_in_28_AWLOCK),
    .m_axi_AWPROT(m_axi_in_28_AWPROT),
    .m_axi_AWQOS(m_axi_in_28_AWQOS),
    .m_axi_AWREADY(m_axi_in_28_AWREADY),
    .m_axi_AWSIZE(m_axi_in_28_AWSIZE),
    .m_axi_AWVALID(m_axi_in_28_AWVALID),
    .m_axi_BID(m_axi_in_28_BID),
    .m_axi_BREADY(m_axi_in_28_BREADY),
    .m_axi_BRESP(m_axi_in_28_BRESP),
    .m_axi_BVALID(m_axi_in_28_BVALID),
    .m_axi_RDATA(m_axi_in_28_RDATA),
    .m_axi_RID(m_axi_in_28_RID),
    .m_axi_RLAST(m_axi_in_28_RLAST),
    .m_axi_RREADY(m_axi_in_28_RREADY),
    .m_axi_RRESP(m_axi_in_28_RRESP),
    .m_axi_RVALID(m_axi_in_28_RVALID),
    .m_axi_WDATA(m_axi_in_28_WDATA),
    .m_axi_WLAST(m_axi_in_28_WLAST),
    .m_axi_WREADY(m_axi_in_28_WREADY),
    .m_axi_WSTRB(m_axi_in_28_WSTRB),
    .m_axi_WVALID(m_axi_in_28_WVALID),
    .read_addr_din(in_28_read_addr__din),
    .read_addr_full_n(in_28_read_addr__full_n),
    .read_addr_write(in_28_read_addr__write),
    .read_data_dout(in_28_read_data__dout),
    .read_data_empty_n(in_28_read_data__empty_n),
    .read_data_read(in_28_read_data__read),
    .write_addr_din(in_28_write_addr__din),
    .write_addr_full_n(in_28_write_addr__full_n),
    .write_addr_write(in_28_write_addr__write),
    .write_data_din(in_28_write_data__din),
    .write_data_full_n(in_28_write_data__full_n),
    .write_data_write(in_28_write_data__write),
    .write_resp_dout(in_28_write_resp__dout),
    .write_resp_empty_n(in_28_write_resp__empty_n),
    .write_resp_read(in_28_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_29__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_29_ARADDR),
    .m_axi_ARBURST(m_axi_in_29_ARBURST),
    .m_axi_ARCACHE(m_axi_in_29_ARCACHE),
    .m_axi_ARID(m_axi_in_29_ARID),
    .m_axi_ARLEN(m_axi_in_29_ARLEN),
    .m_axi_ARLOCK(m_axi_in_29_ARLOCK),
    .m_axi_ARPROT(m_axi_in_29_ARPROT),
    .m_axi_ARQOS(m_axi_in_29_ARQOS),
    .m_axi_ARREADY(m_axi_in_29_ARREADY),
    .m_axi_ARSIZE(m_axi_in_29_ARSIZE),
    .m_axi_ARVALID(m_axi_in_29_ARVALID),
    .m_axi_AWADDR(m_axi_in_29_AWADDR),
    .m_axi_AWBURST(m_axi_in_29_AWBURST),
    .m_axi_AWCACHE(m_axi_in_29_AWCACHE),
    .m_axi_AWID(m_axi_in_29_AWID),
    .m_axi_AWLEN(m_axi_in_29_AWLEN),
    .m_axi_AWLOCK(m_axi_in_29_AWLOCK),
    .m_axi_AWPROT(m_axi_in_29_AWPROT),
    .m_axi_AWQOS(m_axi_in_29_AWQOS),
    .m_axi_AWREADY(m_axi_in_29_AWREADY),
    .m_axi_AWSIZE(m_axi_in_29_AWSIZE),
    .m_axi_AWVALID(m_axi_in_29_AWVALID),
    .m_axi_BID(m_axi_in_29_BID),
    .m_axi_BREADY(m_axi_in_29_BREADY),
    .m_axi_BRESP(m_axi_in_29_BRESP),
    .m_axi_BVALID(m_axi_in_29_BVALID),
    .m_axi_RDATA(m_axi_in_29_RDATA),
    .m_axi_RID(m_axi_in_29_RID),
    .m_axi_RLAST(m_axi_in_29_RLAST),
    .m_axi_RREADY(m_axi_in_29_RREADY),
    .m_axi_RRESP(m_axi_in_29_RRESP),
    .m_axi_RVALID(m_axi_in_29_RVALID),
    .m_axi_WDATA(m_axi_in_29_WDATA),
    .m_axi_WLAST(m_axi_in_29_WLAST),
    .m_axi_WREADY(m_axi_in_29_WREADY),
    .m_axi_WSTRB(m_axi_in_29_WSTRB),
    .m_axi_WVALID(m_axi_in_29_WVALID),
    .read_addr_din(in_29_read_addr__din),
    .read_addr_full_n(in_29_read_addr__full_n),
    .read_addr_write(in_29_read_addr__write),
    .read_data_dout(in_29_read_data__dout),
    .read_data_empty_n(in_29_read_data__empty_n),
    .read_data_read(in_29_read_data__read),
    .write_addr_din(in_29_write_addr__din),
    .write_addr_full_n(in_29_write_addr__full_n),
    .write_addr_write(in_29_write_addr__write),
    .write_data_din(in_29_write_data__din),
    .write_data_full_n(in_29_write_data__full_n),
    .write_data_write(in_29_write_data__write),
    .write_resp_dout(in_29_write_resp__dout),
    .write_resp_empty_n(in_29_write_resp__empty_n),
    .write_resp_read(in_29_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_3_ARADDR),
    .m_axi_ARBURST(m_axi_in_3_ARBURST),
    .m_axi_ARCACHE(m_axi_in_3_ARCACHE),
    .m_axi_ARID(m_axi_in_3_ARID),
    .m_axi_ARLEN(m_axi_in_3_ARLEN),
    .m_axi_ARLOCK(m_axi_in_3_ARLOCK),
    .m_axi_ARPROT(m_axi_in_3_ARPROT),
    .m_axi_ARQOS(m_axi_in_3_ARQOS),
    .m_axi_ARREADY(m_axi_in_3_ARREADY),
    .m_axi_ARSIZE(m_axi_in_3_ARSIZE),
    .m_axi_ARVALID(m_axi_in_3_ARVALID),
    .m_axi_AWADDR(m_axi_in_3_AWADDR),
    .m_axi_AWBURST(m_axi_in_3_AWBURST),
    .m_axi_AWCACHE(m_axi_in_3_AWCACHE),
    .m_axi_AWID(m_axi_in_3_AWID),
    .m_axi_AWLEN(m_axi_in_3_AWLEN),
    .m_axi_AWLOCK(m_axi_in_3_AWLOCK),
    .m_axi_AWPROT(m_axi_in_3_AWPROT),
    .m_axi_AWQOS(m_axi_in_3_AWQOS),
    .m_axi_AWREADY(m_axi_in_3_AWREADY),
    .m_axi_AWSIZE(m_axi_in_3_AWSIZE),
    .m_axi_AWVALID(m_axi_in_3_AWVALID),
    .m_axi_BID(m_axi_in_3_BID),
    .m_axi_BREADY(m_axi_in_3_BREADY),
    .m_axi_BRESP(m_axi_in_3_BRESP),
    .m_axi_BVALID(m_axi_in_3_BVALID),
    .m_axi_RDATA(m_axi_in_3_RDATA),
    .m_axi_RID(m_axi_in_3_RID),
    .m_axi_RLAST(m_axi_in_3_RLAST),
    .m_axi_RREADY(m_axi_in_3_RREADY),
    .m_axi_RRESP(m_axi_in_3_RRESP),
    .m_axi_RVALID(m_axi_in_3_RVALID),
    .m_axi_WDATA(m_axi_in_3_WDATA),
    .m_axi_WLAST(m_axi_in_3_WLAST),
    .m_axi_WREADY(m_axi_in_3_WREADY),
    .m_axi_WSTRB(m_axi_in_3_WSTRB),
    .m_axi_WVALID(m_axi_in_3_WVALID),
    .read_addr_din(in_3_read_addr__din),
    .read_addr_full_n(in_3_read_addr__full_n),
    .read_addr_write(in_3_read_addr__write),
    .read_data_dout(in_3_read_data__dout),
    .read_data_empty_n(in_3_read_data__empty_n),
    .read_data_read(in_3_read_data__read),
    .write_addr_din(in_3_write_addr__din),
    .write_addr_full_n(in_3_write_addr__full_n),
    .write_addr_write(in_3_write_addr__write),
    .write_data_din(in_3_write_data__din),
    .write_data_full_n(in_3_write_data__full_n),
    .write_data_write(in_3_write_data__write),
    .write_resp_dout(in_3_write_resp__dout),
    .write_resp_empty_n(in_3_write_resp__empty_n),
    .write_resp_read(in_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_30__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_30_ARADDR),
    .m_axi_ARBURST(m_axi_in_30_ARBURST),
    .m_axi_ARCACHE(m_axi_in_30_ARCACHE),
    .m_axi_ARID(m_axi_in_30_ARID),
    .m_axi_ARLEN(m_axi_in_30_ARLEN),
    .m_axi_ARLOCK(m_axi_in_30_ARLOCK),
    .m_axi_ARPROT(m_axi_in_30_ARPROT),
    .m_axi_ARQOS(m_axi_in_30_ARQOS),
    .m_axi_ARREADY(m_axi_in_30_ARREADY),
    .m_axi_ARSIZE(m_axi_in_30_ARSIZE),
    .m_axi_ARVALID(m_axi_in_30_ARVALID),
    .m_axi_AWADDR(m_axi_in_30_AWADDR),
    .m_axi_AWBURST(m_axi_in_30_AWBURST),
    .m_axi_AWCACHE(m_axi_in_30_AWCACHE),
    .m_axi_AWID(m_axi_in_30_AWID),
    .m_axi_AWLEN(m_axi_in_30_AWLEN),
    .m_axi_AWLOCK(m_axi_in_30_AWLOCK),
    .m_axi_AWPROT(m_axi_in_30_AWPROT),
    .m_axi_AWQOS(m_axi_in_30_AWQOS),
    .m_axi_AWREADY(m_axi_in_30_AWREADY),
    .m_axi_AWSIZE(m_axi_in_30_AWSIZE),
    .m_axi_AWVALID(m_axi_in_30_AWVALID),
    .m_axi_BID(m_axi_in_30_BID),
    .m_axi_BREADY(m_axi_in_30_BREADY),
    .m_axi_BRESP(m_axi_in_30_BRESP),
    .m_axi_BVALID(m_axi_in_30_BVALID),
    .m_axi_RDATA(m_axi_in_30_RDATA),
    .m_axi_RID(m_axi_in_30_RID),
    .m_axi_RLAST(m_axi_in_30_RLAST),
    .m_axi_RREADY(m_axi_in_30_RREADY),
    .m_axi_RRESP(m_axi_in_30_RRESP),
    .m_axi_RVALID(m_axi_in_30_RVALID),
    .m_axi_WDATA(m_axi_in_30_WDATA),
    .m_axi_WLAST(m_axi_in_30_WLAST),
    .m_axi_WREADY(m_axi_in_30_WREADY),
    .m_axi_WSTRB(m_axi_in_30_WSTRB),
    .m_axi_WVALID(m_axi_in_30_WVALID),
    .read_addr_din(in_30_read_addr__din),
    .read_addr_full_n(in_30_read_addr__full_n),
    .read_addr_write(in_30_read_addr__write),
    .read_data_dout(in_30_read_data__dout),
    .read_data_empty_n(in_30_read_data__empty_n),
    .read_data_read(in_30_read_data__read),
    .write_addr_din(in_30_write_addr__din),
    .write_addr_full_n(in_30_write_addr__full_n),
    .write_addr_write(in_30_write_addr__write),
    .write_data_din(in_30_write_data__din),
    .write_data_full_n(in_30_write_data__full_n),
    .write_data_write(in_30_write_data__write),
    .write_resp_dout(in_30_write_resp__dout),
    .write_resp_empty_n(in_30_write_resp__empty_n),
    .write_resp_read(in_30_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_31__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_31_ARADDR),
    .m_axi_ARBURST(m_axi_in_31_ARBURST),
    .m_axi_ARCACHE(m_axi_in_31_ARCACHE),
    .m_axi_ARID(m_axi_in_31_ARID),
    .m_axi_ARLEN(m_axi_in_31_ARLEN),
    .m_axi_ARLOCK(m_axi_in_31_ARLOCK),
    .m_axi_ARPROT(m_axi_in_31_ARPROT),
    .m_axi_ARQOS(m_axi_in_31_ARQOS),
    .m_axi_ARREADY(m_axi_in_31_ARREADY),
    .m_axi_ARSIZE(m_axi_in_31_ARSIZE),
    .m_axi_ARVALID(m_axi_in_31_ARVALID),
    .m_axi_AWADDR(m_axi_in_31_AWADDR),
    .m_axi_AWBURST(m_axi_in_31_AWBURST),
    .m_axi_AWCACHE(m_axi_in_31_AWCACHE),
    .m_axi_AWID(m_axi_in_31_AWID),
    .m_axi_AWLEN(m_axi_in_31_AWLEN),
    .m_axi_AWLOCK(m_axi_in_31_AWLOCK),
    .m_axi_AWPROT(m_axi_in_31_AWPROT),
    .m_axi_AWQOS(m_axi_in_31_AWQOS),
    .m_axi_AWREADY(m_axi_in_31_AWREADY),
    .m_axi_AWSIZE(m_axi_in_31_AWSIZE),
    .m_axi_AWVALID(m_axi_in_31_AWVALID),
    .m_axi_BID(m_axi_in_31_BID),
    .m_axi_BREADY(m_axi_in_31_BREADY),
    .m_axi_BRESP(m_axi_in_31_BRESP),
    .m_axi_BVALID(m_axi_in_31_BVALID),
    .m_axi_RDATA(m_axi_in_31_RDATA),
    .m_axi_RID(m_axi_in_31_RID),
    .m_axi_RLAST(m_axi_in_31_RLAST),
    .m_axi_RREADY(m_axi_in_31_RREADY),
    .m_axi_RRESP(m_axi_in_31_RRESP),
    .m_axi_RVALID(m_axi_in_31_RVALID),
    .m_axi_WDATA(m_axi_in_31_WDATA),
    .m_axi_WLAST(m_axi_in_31_WLAST),
    .m_axi_WREADY(m_axi_in_31_WREADY),
    .m_axi_WSTRB(m_axi_in_31_WSTRB),
    .m_axi_WVALID(m_axi_in_31_WVALID),
    .read_addr_din(in_31_read_addr__din),
    .read_addr_full_n(in_31_read_addr__full_n),
    .read_addr_write(in_31_read_addr__write),
    .read_data_dout(in_31_read_data__dout),
    .read_data_empty_n(in_31_read_data__empty_n),
    .read_data_read(in_31_read_data__read),
    .write_addr_din(in_31_write_addr__din),
    .write_addr_full_n(in_31_write_addr__full_n),
    .write_addr_write(in_31_write_addr__write),
    .write_data_din(in_31_write_data__din),
    .write_data_full_n(in_31_write_data__full_n),
    .write_data_write(in_31_write_data__write),
    .write_resp_dout(in_31_write_resp__dout),
    .write_resp_empty_n(in_31_write_resp__empty_n),
    .write_resp_read(in_31_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_32__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_32_ARADDR),
    .m_axi_ARBURST(m_axi_in_32_ARBURST),
    .m_axi_ARCACHE(m_axi_in_32_ARCACHE),
    .m_axi_ARID(m_axi_in_32_ARID),
    .m_axi_ARLEN(m_axi_in_32_ARLEN),
    .m_axi_ARLOCK(m_axi_in_32_ARLOCK),
    .m_axi_ARPROT(m_axi_in_32_ARPROT),
    .m_axi_ARQOS(m_axi_in_32_ARQOS),
    .m_axi_ARREADY(m_axi_in_32_ARREADY),
    .m_axi_ARSIZE(m_axi_in_32_ARSIZE),
    .m_axi_ARVALID(m_axi_in_32_ARVALID),
    .m_axi_AWADDR(m_axi_in_32_AWADDR),
    .m_axi_AWBURST(m_axi_in_32_AWBURST),
    .m_axi_AWCACHE(m_axi_in_32_AWCACHE),
    .m_axi_AWID(m_axi_in_32_AWID),
    .m_axi_AWLEN(m_axi_in_32_AWLEN),
    .m_axi_AWLOCK(m_axi_in_32_AWLOCK),
    .m_axi_AWPROT(m_axi_in_32_AWPROT),
    .m_axi_AWQOS(m_axi_in_32_AWQOS),
    .m_axi_AWREADY(m_axi_in_32_AWREADY),
    .m_axi_AWSIZE(m_axi_in_32_AWSIZE),
    .m_axi_AWVALID(m_axi_in_32_AWVALID),
    .m_axi_BID(m_axi_in_32_BID),
    .m_axi_BREADY(m_axi_in_32_BREADY),
    .m_axi_BRESP(m_axi_in_32_BRESP),
    .m_axi_BVALID(m_axi_in_32_BVALID),
    .m_axi_RDATA(m_axi_in_32_RDATA),
    .m_axi_RID(m_axi_in_32_RID),
    .m_axi_RLAST(m_axi_in_32_RLAST),
    .m_axi_RREADY(m_axi_in_32_RREADY),
    .m_axi_RRESP(m_axi_in_32_RRESP),
    .m_axi_RVALID(m_axi_in_32_RVALID),
    .m_axi_WDATA(m_axi_in_32_WDATA),
    .m_axi_WLAST(m_axi_in_32_WLAST),
    .m_axi_WREADY(m_axi_in_32_WREADY),
    .m_axi_WSTRB(m_axi_in_32_WSTRB),
    .m_axi_WVALID(m_axi_in_32_WVALID),
    .read_addr_din(in_32_read_addr__din),
    .read_addr_full_n(in_32_read_addr__full_n),
    .read_addr_write(in_32_read_addr__write),
    .read_data_dout(in_32_read_data__dout),
    .read_data_empty_n(in_32_read_data__empty_n),
    .read_data_read(in_32_read_data__read),
    .write_addr_din(in_32_write_addr__din),
    .write_addr_full_n(in_32_write_addr__full_n),
    .write_addr_write(in_32_write_addr__write),
    .write_data_din(in_32_write_data__din),
    .write_data_full_n(in_32_write_data__full_n),
    .write_data_write(in_32_write_data__write),
    .write_resp_dout(in_32_write_resp__dout),
    .write_resp_empty_n(in_32_write_resp__empty_n),
    .write_resp_read(in_32_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_33__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_33_ARADDR),
    .m_axi_ARBURST(m_axi_in_33_ARBURST),
    .m_axi_ARCACHE(m_axi_in_33_ARCACHE),
    .m_axi_ARID(m_axi_in_33_ARID),
    .m_axi_ARLEN(m_axi_in_33_ARLEN),
    .m_axi_ARLOCK(m_axi_in_33_ARLOCK),
    .m_axi_ARPROT(m_axi_in_33_ARPROT),
    .m_axi_ARQOS(m_axi_in_33_ARQOS),
    .m_axi_ARREADY(m_axi_in_33_ARREADY),
    .m_axi_ARSIZE(m_axi_in_33_ARSIZE),
    .m_axi_ARVALID(m_axi_in_33_ARVALID),
    .m_axi_AWADDR(m_axi_in_33_AWADDR),
    .m_axi_AWBURST(m_axi_in_33_AWBURST),
    .m_axi_AWCACHE(m_axi_in_33_AWCACHE),
    .m_axi_AWID(m_axi_in_33_AWID),
    .m_axi_AWLEN(m_axi_in_33_AWLEN),
    .m_axi_AWLOCK(m_axi_in_33_AWLOCK),
    .m_axi_AWPROT(m_axi_in_33_AWPROT),
    .m_axi_AWQOS(m_axi_in_33_AWQOS),
    .m_axi_AWREADY(m_axi_in_33_AWREADY),
    .m_axi_AWSIZE(m_axi_in_33_AWSIZE),
    .m_axi_AWVALID(m_axi_in_33_AWVALID),
    .m_axi_BID(m_axi_in_33_BID),
    .m_axi_BREADY(m_axi_in_33_BREADY),
    .m_axi_BRESP(m_axi_in_33_BRESP),
    .m_axi_BVALID(m_axi_in_33_BVALID),
    .m_axi_RDATA(m_axi_in_33_RDATA),
    .m_axi_RID(m_axi_in_33_RID),
    .m_axi_RLAST(m_axi_in_33_RLAST),
    .m_axi_RREADY(m_axi_in_33_RREADY),
    .m_axi_RRESP(m_axi_in_33_RRESP),
    .m_axi_RVALID(m_axi_in_33_RVALID),
    .m_axi_WDATA(m_axi_in_33_WDATA),
    .m_axi_WLAST(m_axi_in_33_WLAST),
    .m_axi_WREADY(m_axi_in_33_WREADY),
    .m_axi_WSTRB(m_axi_in_33_WSTRB),
    .m_axi_WVALID(m_axi_in_33_WVALID),
    .read_addr_din(in_33_read_addr__din),
    .read_addr_full_n(in_33_read_addr__full_n),
    .read_addr_write(in_33_read_addr__write),
    .read_data_dout(in_33_read_data__dout),
    .read_data_empty_n(in_33_read_data__empty_n),
    .read_data_read(in_33_read_data__read),
    .write_addr_din(in_33_write_addr__din),
    .write_addr_full_n(in_33_write_addr__full_n),
    .write_addr_write(in_33_write_addr__write),
    .write_data_din(in_33_write_data__din),
    .write_data_full_n(in_33_write_data__full_n),
    .write_data_write(in_33_write_data__write),
    .write_resp_dout(in_33_write_resp__dout),
    .write_resp_empty_n(in_33_write_resp__empty_n),
    .write_resp_read(in_33_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_34__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_34_ARADDR),
    .m_axi_ARBURST(m_axi_in_34_ARBURST),
    .m_axi_ARCACHE(m_axi_in_34_ARCACHE),
    .m_axi_ARID(m_axi_in_34_ARID),
    .m_axi_ARLEN(m_axi_in_34_ARLEN),
    .m_axi_ARLOCK(m_axi_in_34_ARLOCK),
    .m_axi_ARPROT(m_axi_in_34_ARPROT),
    .m_axi_ARQOS(m_axi_in_34_ARQOS),
    .m_axi_ARREADY(m_axi_in_34_ARREADY),
    .m_axi_ARSIZE(m_axi_in_34_ARSIZE),
    .m_axi_ARVALID(m_axi_in_34_ARVALID),
    .m_axi_AWADDR(m_axi_in_34_AWADDR),
    .m_axi_AWBURST(m_axi_in_34_AWBURST),
    .m_axi_AWCACHE(m_axi_in_34_AWCACHE),
    .m_axi_AWID(m_axi_in_34_AWID),
    .m_axi_AWLEN(m_axi_in_34_AWLEN),
    .m_axi_AWLOCK(m_axi_in_34_AWLOCK),
    .m_axi_AWPROT(m_axi_in_34_AWPROT),
    .m_axi_AWQOS(m_axi_in_34_AWQOS),
    .m_axi_AWREADY(m_axi_in_34_AWREADY),
    .m_axi_AWSIZE(m_axi_in_34_AWSIZE),
    .m_axi_AWVALID(m_axi_in_34_AWVALID),
    .m_axi_BID(m_axi_in_34_BID),
    .m_axi_BREADY(m_axi_in_34_BREADY),
    .m_axi_BRESP(m_axi_in_34_BRESP),
    .m_axi_BVALID(m_axi_in_34_BVALID),
    .m_axi_RDATA(m_axi_in_34_RDATA),
    .m_axi_RID(m_axi_in_34_RID),
    .m_axi_RLAST(m_axi_in_34_RLAST),
    .m_axi_RREADY(m_axi_in_34_RREADY),
    .m_axi_RRESP(m_axi_in_34_RRESP),
    .m_axi_RVALID(m_axi_in_34_RVALID),
    .m_axi_WDATA(m_axi_in_34_WDATA),
    .m_axi_WLAST(m_axi_in_34_WLAST),
    .m_axi_WREADY(m_axi_in_34_WREADY),
    .m_axi_WSTRB(m_axi_in_34_WSTRB),
    .m_axi_WVALID(m_axi_in_34_WVALID),
    .read_addr_din(in_34_read_addr__din),
    .read_addr_full_n(in_34_read_addr__full_n),
    .read_addr_write(in_34_read_addr__write),
    .read_data_dout(in_34_read_data__dout),
    .read_data_empty_n(in_34_read_data__empty_n),
    .read_data_read(in_34_read_data__read),
    .write_addr_din(in_34_write_addr__din),
    .write_addr_full_n(in_34_write_addr__full_n),
    .write_addr_write(in_34_write_addr__write),
    .write_data_din(in_34_write_data__din),
    .write_data_full_n(in_34_write_data__full_n),
    .write_data_write(in_34_write_data__write),
    .write_resp_dout(in_34_write_resp__dout),
    .write_resp_empty_n(in_34_write_resp__empty_n),
    .write_resp_read(in_34_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_35__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_35_ARADDR),
    .m_axi_ARBURST(m_axi_in_35_ARBURST),
    .m_axi_ARCACHE(m_axi_in_35_ARCACHE),
    .m_axi_ARID(m_axi_in_35_ARID),
    .m_axi_ARLEN(m_axi_in_35_ARLEN),
    .m_axi_ARLOCK(m_axi_in_35_ARLOCK),
    .m_axi_ARPROT(m_axi_in_35_ARPROT),
    .m_axi_ARQOS(m_axi_in_35_ARQOS),
    .m_axi_ARREADY(m_axi_in_35_ARREADY),
    .m_axi_ARSIZE(m_axi_in_35_ARSIZE),
    .m_axi_ARVALID(m_axi_in_35_ARVALID),
    .m_axi_AWADDR(m_axi_in_35_AWADDR),
    .m_axi_AWBURST(m_axi_in_35_AWBURST),
    .m_axi_AWCACHE(m_axi_in_35_AWCACHE),
    .m_axi_AWID(m_axi_in_35_AWID),
    .m_axi_AWLEN(m_axi_in_35_AWLEN),
    .m_axi_AWLOCK(m_axi_in_35_AWLOCK),
    .m_axi_AWPROT(m_axi_in_35_AWPROT),
    .m_axi_AWQOS(m_axi_in_35_AWQOS),
    .m_axi_AWREADY(m_axi_in_35_AWREADY),
    .m_axi_AWSIZE(m_axi_in_35_AWSIZE),
    .m_axi_AWVALID(m_axi_in_35_AWVALID),
    .m_axi_BID(m_axi_in_35_BID),
    .m_axi_BREADY(m_axi_in_35_BREADY),
    .m_axi_BRESP(m_axi_in_35_BRESP),
    .m_axi_BVALID(m_axi_in_35_BVALID),
    .m_axi_RDATA(m_axi_in_35_RDATA),
    .m_axi_RID(m_axi_in_35_RID),
    .m_axi_RLAST(m_axi_in_35_RLAST),
    .m_axi_RREADY(m_axi_in_35_RREADY),
    .m_axi_RRESP(m_axi_in_35_RRESP),
    .m_axi_RVALID(m_axi_in_35_RVALID),
    .m_axi_WDATA(m_axi_in_35_WDATA),
    .m_axi_WLAST(m_axi_in_35_WLAST),
    .m_axi_WREADY(m_axi_in_35_WREADY),
    .m_axi_WSTRB(m_axi_in_35_WSTRB),
    .m_axi_WVALID(m_axi_in_35_WVALID),
    .read_addr_din(in_35_read_addr__din),
    .read_addr_full_n(in_35_read_addr__full_n),
    .read_addr_write(in_35_read_addr__write),
    .read_data_dout(in_35_read_data__dout),
    .read_data_empty_n(in_35_read_data__empty_n),
    .read_data_read(in_35_read_data__read),
    .write_addr_din(in_35_write_addr__din),
    .write_addr_full_n(in_35_write_addr__full_n),
    .write_addr_write(in_35_write_addr__write),
    .write_data_din(in_35_write_data__din),
    .write_data_full_n(in_35_write_data__full_n),
    .write_data_write(in_35_write_data__write),
    .write_resp_dout(in_35_write_resp__dout),
    .write_resp_empty_n(in_35_write_resp__empty_n),
    .write_resp_read(in_35_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_36__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_36_ARADDR),
    .m_axi_ARBURST(m_axi_in_36_ARBURST),
    .m_axi_ARCACHE(m_axi_in_36_ARCACHE),
    .m_axi_ARID(m_axi_in_36_ARID),
    .m_axi_ARLEN(m_axi_in_36_ARLEN),
    .m_axi_ARLOCK(m_axi_in_36_ARLOCK),
    .m_axi_ARPROT(m_axi_in_36_ARPROT),
    .m_axi_ARQOS(m_axi_in_36_ARQOS),
    .m_axi_ARREADY(m_axi_in_36_ARREADY),
    .m_axi_ARSIZE(m_axi_in_36_ARSIZE),
    .m_axi_ARVALID(m_axi_in_36_ARVALID),
    .m_axi_AWADDR(m_axi_in_36_AWADDR),
    .m_axi_AWBURST(m_axi_in_36_AWBURST),
    .m_axi_AWCACHE(m_axi_in_36_AWCACHE),
    .m_axi_AWID(m_axi_in_36_AWID),
    .m_axi_AWLEN(m_axi_in_36_AWLEN),
    .m_axi_AWLOCK(m_axi_in_36_AWLOCK),
    .m_axi_AWPROT(m_axi_in_36_AWPROT),
    .m_axi_AWQOS(m_axi_in_36_AWQOS),
    .m_axi_AWREADY(m_axi_in_36_AWREADY),
    .m_axi_AWSIZE(m_axi_in_36_AWSIZE),
    .m_axi_AWVALID(m_axi_in_36_AWVALID),
    .m_axi_BID(m_axi_in_36_BID),
    .m_axi_BREADY(m_axi_in_36_BREADY),
    .m_axi_BRESP(m_axi_in_36_BRESP),
    .m_axi_BVALID(m_axi_in_36_BVALID),
    .m_axi_RDATA(m_axi_in_36_RDATA),
    .m_axi_RID(m_axi_in_36_RID),
    .m_axi_RLAST(m_axi_in_36_RLAST),
    .m_axi_RREADY(m_axi_in_36_RREADY),
    .m_axi_RRESP(m_axi_in_36_RRESP),
    .m_axi_RVALID(m_axi_in_36_RVALID),
    .m_axi_WDATA(m_axi_in_36_WDATA),
    .m_axi_WLAST(m_axi_in_36_WLAST),
    .m_axi_WREADY(m_axi_in_36_WREADY),
    .m_axi_WSTRB(m_axi_in_36_WSTRB),
    .m_axi_WVALID(m_axi_in_36_WVALID),
    .read_addr_din(in_36_read_addr__din),
    .read_addr_full_n(in_36_read_addr__full_n),
    .read_addr_write(in_36_read_addr__write),
    .read_data_dout(in_36_read_data__dout),
    .read_data_empty_n(in_36_read_data__empty_n),
    .read_data_read(in_36_read_data__read),
    .write_addr_din(in_36_write_addr__din),
    .write_addr_full_n(in_36_write_addr__full_n),
    .write_addr_write(in_36_write_addr__write),
    .write_data_din(in_36_write_data__din),
    .write_data_full_n(in_36_write_data__full_n),
    .write_data_write(in_36_write_data__write),
    .write_resp_dout(in_36_write_resp__dout),
    .write_resp_empty_n(in_36_write_resp__empty_n),
    .write_resp_read(in_36_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_37__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_37_ARADDR),
    .m_axi_ARBURST(m_axi_in_37_ARBURST),
    .m_axi_ARCACHE(m_axi_in_37_ARCACHE),
    .m_axi_ARID(m_axi_in_37_ARID),
    .m_axi_ARLEN(m_axi_in_37_ARLEN),
    .m_axi_ARLOCK(m_axi_in_37_ARLOCK),
    .m_axi_ARPROT(m_axi_in_37_ARPROT),
    .m_axi_ARQOS(m_axi_in_37_ARQOS),
    .m_axi_ARREADY(m_axi_in_37_ARREADY),
    .m_axi_ARSIZE(m_axi_in_37_ARSIZE),
    .m_axi_ARVALID(m_axi_in_37_ARVALID),
    .m_axi_AWADDR(m_axi_in_37_AWADDR),
    .m_axi_AWBURST(m_axi_in_37_AWBURST),
    .m_axi_AWCACHE(m_axi_in_37_AWCACHE),
    .m_axi_AWID(m_axi_in_37_AWID),
    .m_axi_AWLEN(m_axi_in_37_AWLEN),
    .m_axi_AWLOCK(m_axi_in_37_AWLOCK),
    .m_axi_AWPROT(m_axi_in_37_AWPROT),
    .m_axi_AWQOS(m_axi_in_37_AWQOS),
    .m_axi_AWREADY(m_axi_in_37_AWREADY),
    .m_axi_AWSIZE(m_axi_in_37_AWSIZE),
    .m_axi_AWVALID(m_axi_in_37_AWVALID),
    .m_axi_BID(m_axi_in_37_BID),
    .m_axi_BREADY(m_axi_in_37_BREADY),
    .m_axi_BRESP(m_axi_in_37_BRESP),
    .m_axi_BVALID(m_axi_in_37_BVALID),
    .m_axi_RDATA(m_axi_in_37_RDATA),
    .m_axi_RID(m_axi_in_37_RID),
    .m_axi_RLAST(m_axi_in_37_RLAST),
    .m_axi_RREADY(m_axi_in_37_RREADY),
    .m_axi_RRESP(m_axi_in_37_RRESP),
    .m_axi_RVALID(m_axi_in_37_RVALID),
    .m_axi_WDATA(m_axi_in_37_WDATA),
    .m_axi_WLAST(m_axi_in_37_WLAST),
    .m_axi_WREADY(m_axi_in_37_WREADY),
    .m_axi_WSTRB(m_axi_in_37_WSTRB),
    .m_axi_WVALID(m_axi_in_37_WVALID),
    .read_addr_din(in_37_read_addr__din),
    .read_addr_full_n(in_37_read_addr__full_n),
    .read_addr_write(in_37_read_addr__write),
    .read_data_dout(in_37_read_data__dout),
    .read_data_empty_n(in_37_read_data__empty_n),
    .read_data_read(in_37_read_data__read),
    .write_addr_din(in_37_write_addr__din),
    .write_addr_full_n(in_37_write_addr__full_n),
    .write_addr_write(in_37_write_addr__write),
    .write_data_din(in_37_write_data__din),
    .write_data_full_n(in_37_write_data__full_n),
    .write_data_write(in_37_write_data__write),
    .write_resp_dout(in_37_write_resp__dout),
    .write_resp_empty_n(in_37_write_resp__empty_n),
    .write_resp_read(in_37_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_38__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_38_ARADDR),
    .m_axi_ARBURST(m_axi_in_38_ARBURST),
    .m_axi_ARCACHE(m_axi_in_38_ARCACHE),
    .m_axi_ARID(m_axi_in_38_ARID),
    .m_axi_ARLEN(m_axi_in_38_ARLEN),
    .m_axi_ARLOCK(m_axi_in_38_ARLOCK),
    .m_axi_ARPROT(m_axi_in_38_ARPROT),
    .m_axi_ARQOS(m_axi_in_38_ARQOS),
    .m_axi_ARREADY(m_axi_in_38_ARREADY),
    .m_axi_ARSIZE(m_axi_in_38_ARSIZE),
    .m_axi_ARVALID(m_axi_in_38_ARVALID),
    .m_axi_AWADDR(m_axi_in_38_AWADDR),
    .m_axi_AWBURST(m_axi_in_38_AWBURST),
    .m_axi_AWCACHE(m_axi_in_38_AWCACHE),
    .m_axi_AWID(m_axi_in_38_AWID),
    .m_axi_AWLEN(m_axi_in_38_AWLEN),
    .m_axi_AWLOCK(m_axi_in_38_AWLOCK),
    .m_axi_AWPROT(m_axi_in_38_AWPROT),
    .m_axi_AWQOS(m_axi_in_38_AWQOS),
    .m_axi_AWREADY(m_axi_in_38_AWREADY),
    .m_axi_AWSIZE(m_axi_in_38_AWSIZE),
    .m_axi_AWVALID(m_axi_in_38_AWVALID),
    .m_axi_BID(m_axi_in_38_BID),
    .m_axi_BREADY(m_axi_in_38_BREADY),
    .m_axi_BRESP(m_axi_in_38_BRESP),
    .m_axi_BVALID(m_axi_in_38_BVALID),
    .m_axi_RDATA(m_axi_in_38_RDATA),
    .m_axi_RID(m_axi_in_38_RID),
    .m_axi_RLAST(m_axi_in_38_RLAST),
    .m_axi_RREADY(m_axi_in_38_RREADY),
    .m_axi_RRESP(m_axi_in_38_RRESP),
    .m_axi_RVALID(m_axi_in_38_RVALID),
    .m_axi_WDATA(m_axi_in_38_WDATA),
    .m_axi_WLAST(m_axi_in_38_WLAST),
    .m_axi_WREADY(m_axi_in_38_WREADY),
    .m_axi_WSTRB(m_axi_in_38_WSTRB),
    .m_axi_WVALID(m_axi_in_38_WVALID),
    .read_addr_din(in_38_read_addr__din),
    .read_addr_full_n(in_38_read_addr__full_n),
    .read_addr_write(in_38_read_addr__write),
    .read_data_dout(in_38_read_data__dout),
    .read_data_empty_n(in_38_read_data__empty_n),
    .read_data_read(in_38_read_data__read),
    .write_addr_din(in_38_write_addr__din),
    .write_addr_full_n(in_38_write_addr__full_n),
    .write_addr_write(in_38_write_addr__write),
    .write_data_din(in_38_write_data__din),
    .write_data_full_n(in_38_write_data__full_n),
    .write_data_write(in_38_write_data__write),
    .write_resp_dout(in_38_write_resp__dout),
    .write_resp_empty_n(in_38_write_resp__empty_n),
    .write_resp_read(in_38_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_39__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_39_ARADDR),
    .m_axi_ARBURST(m_axi_in_39_ARBURST),
    .m_axi_ARCACHE(m_axi_in_39_ARCACHE),
    .m_axi_ARID(m_axi_in_39_ARID),
    .m_axi_ARLEN(m_axi_in_39_ARLEN),
    .m_axi_ARLOCK(m_axi_in_39_ARLOCK),
    .m_axi_ARPROT(m_axi_in_39_ARPROT),
    .m_axi_ARQOS(m_axi_in_39_ARQOS),
    .m_axi_ARREADY(m_axi_in_39_ARREADY),
    .m_axi_ARSIZE(m_axi_in_39_ARSIZE),
    .m_axi_ARVALID(m_axi_in_39_ARVALID),
    .m_axi_AWADDR(m_axi_in_39_AWADDR),
    .m_axi_AWBURST(m_axi_in_39_AWBURST),
    .m_axi_AWCACHE(m_axi_in_39_AWCACHE),
    .m_axi_AWID(m_axi_in_39_AWID),
    .m_axi_AWLEN(m_axi_in_39_AWLEN),
    .m_axi_AWLOCK(m_axi_in_39_AWLOCK),
    .m_axi_AWPROT(m_axi_in_39_AWPROT),
    .m_axi_AWQOS(m_axi_in_39_AWQOS),
    .m_axi_AWREADY(m_axi_in_39_AWREADY),
    .m_axi_AWSIZE(m_axi_in_39_AWSIZE),
    .m_axi_AWVALID(m_axi_in_39_AWVALID),
    .m_axi_BID(m_axi_in_39_BID),
    .m_axi_BREADY(m_axi_in_39_BREADY),
    .m_axi_BRESP(m_axi_in_39_BRESP),
    .m_axi_BVALID(m_axi_in_39_BVALID),
    .m_axi_RDATA(m_axi_in_39_RDATA),
    .m_axi_RID(m_axi_in_39_RID),
    .m_axi_RLAST(m_axi_in_39_RLAST),
    .m_axi_RREADY(m_axi_in_39_RREADY),
    .m_axi_RRESP(m_axi_in_39_RRESP),
    .m_axi_RVALID(m_axi_in_39_RVALID),
    .m_axi_WDATA(m_axi_in_39_WDATA),
    .m_axi_WLAST(m_axi_in_39_WLAST),
    .m_axi_WREADY(m_axi_in_39_WREADY),
    .m_axi_WSTRB(m_axi_in_39_WSTRB),
    .m_axi_WVALID(m_axi_in_39_WVALID),
    .read_addr_din(in_39_read_addr__din),
    .read_addr_full_n(in_39_read_addr__full_n),
    .read_addr_write(in_39_read_addr__write),
    .read_data_dout(in_39_read_data__dout),
    .read_data_empty_n(in_39_read_data__empty_n),
    .read_data_read(in_39_read_data__read),
    .write_addr_din(in_39_write_addr__din),
    .write_addr_full_n(in_39_write_addr__full_n),
    .write_addr_write(in_39_write_addr__write),
    .write_data_din(in_39_write_data__din),
    .write_data_full_n(in_39_write_data__full_n),
    .write_data_write(in_39_write_data__write),
    .write_resp_dout(in_39_write_resp__dout),
    .write_resp_empty_n(in_39_write_resp__empty_n),
    .write_resp_read(in_39_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_4_ARADDR),
    .m_axi_ARBURST(m_axi_in_4_ARBURST),
    .m_axi_ARCACHE(m_axi_in_4_ARCACHE),
    .m_axi_ARID(m_axi_in_4_ARID),
    .m_axi_ARLEN(m_axi_in_4_ARLEN),
    .m_axi_ARLOCK(m_axi_in_4_ARLOCK),
    .m_axi_ARPROT(m_axi_in_4_ARPROT),
    .m_axi_ARQOS(m_axi_in_4_ARQOS),
    .m_axi_ARREADY(m_axi_in_4_ARREADY),
    .m_axi_ARSIZE(m_axi_in_4_ARSIZE),
    .m_axi_ARVALID(m_axi_in_4_ARVALID),
    .m_axi_AWADDR(m_axi_in_4_AWADDR),
    .m_axi_AWBURST(m_axi_in_4_AWBURST),
    .m_axi_AWCACHE(m_axi_in_4_AWCACHE),
    .m_axi_AWID(m_axi_in_4_AWID),
    .m_axi_AWLEN(m_axi_in_4_AWLEN),
    .m_axi_AWLOCK(m_axi_in_4_AWLOCK),
    .m_axi_AWPROT(m_axi_in_4_AWPROT),
    .m_axi_AWQOS(m_axi_in_4_AWQOS),
    .m_axi_AWREADY(m_axi_in_4_AWREADY),
    .m_axi_AWSIZE(m_axi_in_4_AWSIZE),
    .m_axi_AWVALID(m_axi_in_4_AWVALID),
    .m_axi_BID(m_axi_in_4_BID),
    .m_axi_BREADY(m_axi_in_4_BREADY),
    .m_axi_BRESP(m_axi_in_4_BRESP),
    .m_axi_BVALID(m_axi_in_4_BVALID),
    .m_axi_RDATA(m_axi_in_4_RDATA),
    .m_axi_RID(m_axi_in_4_RID),
    .m_axi_RLAST(m_axi_in_4_RLAST),
    .m_axi_RREADY(m_axi_in_4_RREADY),
    .m_axi_RRESP(m_axi_in_4_RRESP),
    .m_axi_RVALID(m_axi_in_4_RVALID),
    .m_axi_WDATA(m_axi_in_4_WDATA),
    .m_axi_WLAST(m_axi_in_4_WLAST),
    .m_axi_WREADY(m_axi_in_4_WREADY),
    .m_axi_WSTRB(m_axi_in_4_WSTRB),
    .m_axi_WVALID(m_axi_in_4_WVALID),
    .read_addr_din(in_4_read_addr__din),
    .read_addr_full_n(in_4_read_addr__full_n),
    .read_addr_write(in_4_read_addr__write),
    .read_data_dout(in_4_read_data__dout),
    .read_data_empty_n(in_4_read_data__empty_n),
    .read_data_read(in_4_read_data__read),
    .write_addr_din(in_4_write_addr__din),
    .write_addr_full_n(in_4_write_addr__full_n),
    .write_addr_write(in_4_write_addr__write),
    .write_data_din(in_4_write_data__din),
    .write_data_full_n(in_4_write_data__full_n),
    .write_data_write(in_4_write_data__write),
    .write_resp_dout(in_4_write_resp__dout),
    .write_resp_empty_n(in_4_write_resp__empty_n),
    .write_resp_read(in_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_40__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_40_ARADDR),
    .m_axi_ARBURST(m_axi_in_40_ARBURST),
    .m_axi_ARCACHE(m_axi_in_40_ARCACHE),
    .m_axi_ARID(m_axi_in_40_ARID),
    .m_axi_ARLEN(m_axi_in_40_ARLEN),
    .m_axi_ARLOCK(m_axi_in_40_ARLOCK),
    .m_axi_ARPROT(m_axi_in_40_ARPROT),
    .m_axi_ARQOS(m_axi_in_40_ARQOS),
    .m_axi_ARREADY(m_axi_in_40_ARREADY),
    .m_axi_ARSIZE(m_axi_in_40_ARSIZE),
    .m_axi_ARVALID(m_axi_in_40_ARVALID),
    .m_axi_AWADDR(m_axi_in_40_AWADDR),
    .m_axi_AWBURST(m_axi_in_40_AWBURST),
    .m_axi_AWCACHE(m_axi_in_40_AWCACHE),
    .m_axi_AWID(m_axi_in_40_AWID),
    .m_axi_AWLEN(m_axi_in_40_AWLEN),
    .m_axi_AWLOCK(m_axi_in_40_AWLOCK),
    .m_axi_AWPROT(m_axi_in_40_AWPROT),
    .m_axi_AWQOS(m_axi_in_40_AWQOS),
    .m_axi_AWREADY(m_axi_in_40_AWREADY),
    .m_axi_AWSIZE(m_axi_in_40_AWSIZE),
    .m_axi_AWVALID(m_axi_in_40_AWVALID),
    .m_axi_BID(m_axi_in_40_BID),
    .m_axi_BREADY(m_axi_in_40_BREADY),
    .m_axi_BRESP(m_axi_in_40_BRESP),
    .m_axi_BVALID(m_axi_in_40_BVALID),
    .m_axi_RDATA(m_axi_in_40_RDATA),
    .m_axi_RID(m_axi_in_40_RID),
    .m_axi_RLAST(m_axi_in_40_RLAST),
    .m_axi_RREADY(m_axi_in_40_RREADY),
    .m_axi_RRESP(m_axi_in_40_RRESP),
    .m_axi_RVALID(m_axi_in_40_RVALID),
    .m_axi_WDATA(m_axi_in_40_WDATA),
    .m_axi_WLAST(m_axi_in_40_WLAST),
    .m_axi_WREADY(m_axi_in_40_WREADY),
    .m_axi_WSTRB(m_axi_in_40_WSTRB),
    .m_axi_WVALID(m_axi_in_40_WVALID),
    .read_addr_din(in_40_read_addr__din),
    .read_addr_full_n(in_40_read_addr__full_n),
    .read_addr_write(in_40_read_addr__write),
    .read_data_dout(in_40_read_data__dout),
    .read_data_empty_n(in_40_read_data__empty_n),
    .read_data_read(in_40_read_data__read),
    .write_addr_din(in_40_write_addr__din),
    .write_addr_full_n(in_40_write_addr__full_n),
    .write_addr_write(in_40_write_addr__write),
    .write_data_din(in_40_write_data__din),
    .write_data_full_n(in_40_write_data__full_n),
    .write_data_write(in_40_write_data__write),
    .write_resp_dout(in_40_write_resp__dout),
    .write_resp_empty_n(in_40_write_resp__empty_n),
    .write_resp_read(in_40_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_41__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_41_ARADDR),
    .m_axi_ARBURST(m_axi_in_41_ARBURST),
    .m_axi_ARCACHE(m_axi_in_41_ARCACHE),
    .m_axi_ARID(m_axi_in_41_ARID),
    .m_axi_ARLEN(m_axi_in_41_ARLEN),
    .m_axi_ARLOCK(m_axi_in_41_ARLOCK),
    .m_axi_ARPROT(m_axi_in_41_ARPROT),
    .m_axi_ARQOS(m_axi_in_41_ARQOS),
    .m_axi_ARREADY(m_axi_in_41_ARREADY),
    .m_axi_ARSIZE(m_axi_in_41_ARSIZE),
    .m_axi_ARVALID(m_axi_in_41_ARVALID),
    .m_axi_AWADDR(m_axi_in_41_AWADDR),
    .m_axi_AWBURST(m_axi_in_41_AWBURST),
    .m_axi_AWCACHE(m_axi_in_41_AWCACHE),
    .m_axi_AWID(m_axi_in_41_AWID),
    .m_axi_AWLEN(m_axi_in_41_AWLEN),
    .m_axi_AWLOCK(m_axi_in_41_AWLOCK),
    .m_axi_AWPROT(m_axi_in_41_AWPROT),
    .m_axi_AWQOS(m_axi_in_41_AWQOS),
    .m_axi_AWREADY(m_axi_in_41_AWREADY),
    .m_axi_AWSIZE(m_axi_in_41_AWSIZE),
    .m_axi_AWVALID(m_axi_in_41_AWVALID),
    .m_axi_BID(m_axi_in_41_BID),
    .m_axi_BREADY(m_axi_in_41_BREADY),
    .m_axi_BRESP(m_axi_in_41_BRESP),
    .m_axi_BVALID(m_axi_in_41_BVALID),
    .m_axi_RDATA(m_axi_in_41_RDATA),
    .m_axi_RID(m_axi_in_41_RID),
    .m_axi_RLAST(m_axi_in_41_RLAST),
    .m_axi_RREADY(m_axi_in_41_RREADY),
    .m_axi_RRESP(m_axi_in_41_RRESP),
    .m_axi_RVALID(m_axi_in_41_RVALID),
    .m_axi_WDATA(m_axi_in_41_WDATA),
    .m_axi_WLAST(m_axi_in_41_WLAST),
    .m_axi_WREADY(m_axi_in_41_WREADY),
    .m_axi_WSTRB(m_axi_in_41_WSTRB),
    .m_axi_WVALID(m_axi_in_41_WVALID),
    .read_addr_din(in_41_read_addr__din),
    .read_addr_full_n(in_41_read_addr__full_n),
    .read_addr_write(in_41_read_addr__write),
    .read_data_dout(in_41_read_data__dout),
    .read_data_empty_n(in_41_read_data__empty_n),
    .read_data_read(in_41_read_data__read),
    .write_addr_din(in_41_write_addr__din),
    .write_addr_full_n(in_41_write_addr__full_n),
    .write_addr_write(in_41_write_addr__write),
    .write_data_din(in_41_write_data__din),
    .write_data_full_n(in_41_write_data__full_n),
    .write_data_write(in_41_write_data__write),
    .write_resp_dout(in_41_write_resp__dout),
    .write_resp_empty_n(in_41_write_resp__empty_n),
    .write_resp_read(in_41_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_42__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_42_ARADDR),
    .m_axi_ARBURST(m_axi_in_42_ARBURST),
    .m_axi_ARCACHE(m_axi_in_42_ARCACHE),
    .m_axi_ARID(m_axi_in_42_ARID),
    .m_axi_ARLEN(m_axi_in_42_ARLEN),
    .m_axi_ARLOCK(m_axi_in_42_ARLOCK),
    .m_axi_ARPROT(m_axi_in_42_ARPROT),
    .m_axi_ARQOS(m_axi_in_42_ARQOS),
    .m_axi_ARREADY(m_axi_in_42_ARREADY),
    .m_axi_ARSIZE(m_axi_in_42_ARSIZE),
    .m_axi_ARVALID(m_axi_in_42_ARVALID),
    .m_axi_AWADDR(m_axi_in_42_AWADDR),
    .m_axi_AWBURST(m_axi_in_42_AWBURST),
    .m_axi_AWCACHE(m_axi_in_42_AWCACHE),
    .m_axi_AWID(m_axi_in_42_AWID),
    .m_axi_AWLEN(m_axi_in_42_AWLEN),
    .m_axi_AWLOCK(m_axi_in_42_AWLOCK),
    .m_axi_AWPROT(m_axi_in_42_AWPROT),
    .m_axi_AWQOS(m_axi_in_42_AWQOS),
    .m_axi_AWREADY(m_axi_in_42_AWREADY),
    .m_axi_AWSIZE(m_axi_in_42_AWSIZE),
    .m_axi_AWVALID(m_axi_in_42_AWVALID),
    .m_axi_BID(m_axi_in_42_BID),
    .m_axi_BREADY(m_axi_in_42_BREADY),
    .m_axi_BRESP(m_axi_in_42_BRESP),
    .m_axi_BVALID(m_axi_in_42_BVALID),
    .m_axi_RDATA(m_axi_in_42_RDATA),
    .m_axi_RID(m_axi_in_42_RID),
    .m_axi_RLAST(m_axi_in_42_RLAST),
    .m_axi_RREADY(m_axi_in_42_RREADY),
    .m_axi_RRESP(m_axi_in_42_RRESP),
    .m_axi_RVALID(m_axi_in_42_RVALID),
    .m_axi_WDATA(m_axi_in_42_WDATA),
    .m_axi_WLAST(m_axi_in_42_WLAST),
    .m_axi_WREADY(m_axi_in_42_WREADY),
    .m_axi_WSTRB(m_axi_in_42_WSTRB),
    .m_axi_WVALID(m_axi_in_42_WVALID),
    .read_addr_din(in_42_read_addr__din),
    .read_addr_full_n(in_42_read_addr__full_n),
    .read_addr_write(in_42_read_addr__write),
    .read_data_dout(in_42_read_data__dout),
    .read_data_empty_n(in_42_read_data__empty_n),
    .read_data_read(in_42_read_data__read),
    .write_addr_din(in_42_write_addr__din),
    .write_addr_full_n(in_42_write_addr__full_n),
    .write_addr_write(in_42_write_addr__write),
    .write_data_din(in_42_write_data__din),
    .write_data_full_n(in_42_write_data__full_n),
    .write_data_write(in_42_write_data__write),
    .write_resp_dout(in_42_write_resp__dout),
    .write_resp_empty_n(in_42_write_resp__empty_n),
    .write_resp_read(in_42_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_43__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_43_ARADDR),
    .m_axi_ARBURST(m_axi_in_43_ARBURST),
    .m_axi_ARCACHE(m_axi_in_43_ARCACHE),
    .m_axi_ARID(m_axi_in_43_ARID),
    .m_axi_ARLEN(m_axi_in_43_ARLEN),
    .m_axi_ARLOCK(m_axi_in_43_ARLOCK),
    .m_axi_ARPROT(m_axi_in_43_ARPROT),
    .m_axi_ARQOS(m_axi_in_43_ARQOS),
    .m_axi_ARREADY(m_axi_in_43_ARREADY),
    .m_axi_ARSIZE(m_axi_in_43_ARSIZE),
    .m_axi_ARVALID(m_axi_in_43_ARVALID),
    .m_axi_AWADDR(m_axi_in_43_AWADDR),
    .m_axi_AWBURST(m_axi_in_43_AWBURST),
    .m_axi_AWCACHE(m_axi_in_43_AWCACHE),
    .m_axi_AWID(m_axi_in_43_AWID),
    .m_axi_AWLEN(m_axi_in_43_AWLEN),
    .m_axi_AWLOCK(m_axi_in_43_AWLOCK),
    .m_axi_AWPROT(m_axi_in_43_AWPROT),
    .m_axi_AWQOS(m_axi_in_43_AWQOS),
    .m_axi_AWREADY(m_axi_in_43_AWREADY),
    .m_axi_AWSIZE(m_axi_in_43_AWSIZE),
    .m_axi_AWVALID(m_axi_in_43_AWVALID),
    .m_axi_BID(m_axi_in_43_BID),
    .m_axi_BREADY(m_axi_in_43_BREADY),
    .m_axi_BRESP(m_axi_in_43_BRESP),
    .m_axi_BVALID(m_axi_in_43_BVALID),
    .m_axi_RDATA(m_axi_in_43_RDATA),
    .m_axi_RID(m_axi_in_43_RID),
    .m_axi_RLAST(m_axi_in_43_RLAST),
    .m_axi_RREADY(m_axi_in_43_RREADY),
    .m_axi_RRESP(m_axi_in_43_RRESP),
    .m_axi_RVALID(m_axi_in_43_RVALID),
    .m_axi_WDATA(m_axi_in_43_WDATA),
    .m_axi_WLAST(m_axi_in_43_WLAST),
    .m_axi_WREADY(m_axi_in_43_WREADY),
    .m_axi_WSTRB(m_axi_in_43_WSTRB),
    .m_axi_WVALID(m_axi_in_43_WVALID),
    .read_addr_din(in_43_read_addr__din),
    .read_addr_full_n(in_43_read_addr__full_n),
    .read_addr_write(in_43_read_addr__write),
    .read_data_dout(in_43_read_data__dout),
    .read_data_empty_n(in_43_read_data__empty_n),
    .read_data_read(in_43_read_data__read),
    .write_addr_din(in_43_write_addr__din),
    .write_addr_full_n(in_43_write_addr__full_n),
    .write_addr_write(in_43_write_addr__write),
    .write_data_din(in_43_write_data__din),
    .write_data_full_n(in_43_write_data__full_n),
    .write_data_write(in_43_write_data__write),
    .write_resp_dout(in_43_write_resp__dout),
    .write_resp_empty_n(in_43_write_resp__empty_n),
    .write_resp_read(in_43_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_44__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_44_ARADDR),
    .m_axi_ARBURST(m_axi_in_44_ARBURST),
    .m_axi_ARCACHE(m_axi_in_44_ARCACHE),
    .m_axi_ARID(m_axi_in_44_ARID),
    .m_axi_ARLEN(m_axi_in_44_ARLEN),
    .m_axi_ARLOCK(m_axi_in_44_ARLOCK),
    .m_axi_ARPROT(m_axi_in_44_ARPROT),
    .m_axi_ARQOS(m_axi_in_44_ARQOS),
    .m_axi_ARREADY(m_axi_in_44_ARREADY),
    .m_axi_ARSIZE(m_axi_in_44_ARSIZE),
    .m_axi_ARVALID(m_axi_in_44_ARVALID),
    .m_axi_AWADDR(m_axi_in_44_AWADDR),
    .m_axi_AWBURST(m_axi_in_44_AWBURST),
    .m_axi_AWCACHE(m_axi_in_44_AWCACHE),
    .m_axi_AWID(m_axi_in_44_AWID),
    .m_axi_AWLEN(m_axi_in_44_AWLEN),
    .m_axi_AWLOCK(m_axi_in_44_AWLOCK),
    .m_axi_AWPROT(m_axi_in_44_AWPROT),
    .m_axi_AWQOS(m_axi_in_44_AWQOS),
    .m_axi_AWREADY(m_axi_in_44_AWREADY),
    .m_axi_AWSIZE(m_axi_in_44_AWSIZE),
    .m_axi_AWVALID(m_axi_in_44_AWVALID),
    .m_axi_BID(m_axi_in_44_BID),
    .m_axi_BREADY(m_axi_in_44_BREADY),
    .m_axi_BRESP(m_axi_in_44_BRESP),
    .m_axi_BVALID(m_axi_in_44_BVALID),
    .m_axi_RDATA(m_axi_in_44_RDATA),
    .m_axi_RID(m_axi_in_44_RID),
    .m_axi_RLAST(m_axi_in_44_RLAST),
    .m_axi_RREADY(m_axi_in_44_RREADY),
    .m_axi_RRESP(m_axi_in_44_RRESP),
    .m_axi_RVALID(m_axi_in_44_RVALID),
    .m_axi_WDATA(m_axi_in_44_WDATA),
    .m_axi_WLAST(m_axi_in_44_WLAST),
    .m_axi_WREADY(m_axi_in_44_WREADY),
    .m_axi_WSTRB(m_axi_in_44_WSTRB),
    .m_axi_WVALID(m_axi_in_44_WVALID),
    .read_addr_din(in_44_read_addr__din),
    .read_addr_full_n(in_44_read_addr__full_n),
    .read_addr_write(in_44_read_addr__write),
    .read_data_dout(in_44_read_data__dout),
    .read_data_empty_n(in_44_read_data__empty_n),
    .read_data_read(in_44_read_data__read),
    .write_addr_din(in_44_write_addr__din),
    .write_addr_full_n(in_44_write_addr__full_n),
    .write_addr_write(in_44_write_addr__write),
    .write_data_din(in_44_write_data__din),
    .write_data_full_n(in_44_write_data__full_n),
    .write_data_write(in_44_write_data__write),
    .write_resp_dout(in_44_write_resp__dout),
    .write_resp_empty_n(in_44_write_resp__empty_n),
    .write_resp_read(in_44_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_45__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_45_ARADDR),
    .m_axi_ARBURST(m_axi_in_45_ARBURST),
    .m_axi_ARCACHE(m_axi_in_45_ARCACHE),
    .m_axi_ARID(m_axi_in_45_ARID),
    .m_axi_ARLEN(m_axi_in_45_ARLEN),
    .m_axi_ARLOCK(m_axi_in_45_ARLOCK),
    .m_axi_ARPROT(m_axi_in_45_ARPROT),
    .m_axi_ARQOS(m_axi_in_45_ARQOS),
    .m_axi_ARREADY(m_axi_in_45_ARREADY),
    .m_axi_ARSIZE(m_axi_in_45_ARSIZE),
    .m_axi_ARVALID(m_axi_in_45_ARVALID),
    .m_axi_AWADDR(m_axi_in_45_AWADDR),
    .m_axi_AWBURST(m_axi_in_45_AWBURST),
    .m_axi_AWCACHE(m_axi_in_45_AWCACHE),
    .m_axi_AWID(m_axi_in_45_AWID),
    .m_axi_AWLEN(m_axi_in_45_AWLEN),
    .m_axi_AWLOCK(m_axi_in_45_AWLOCK),
    .m_axi_AWPROT(m_axi_in_45_AWPROT),
    .m_axi_AWQOS(m_axi_in_45_AWQOS),
    .m_axi_AWREADY(m_axi_in_45_AWREADY),
    .m_axi_AWSIZE(m_axi_in_45_AWSIZE),
    .m_axi_AWVALID(m_axi_in_45_AWVALID),
    .m_axi_BID(m_axi_in_45_BID),
    .m_axi_BREADY(m_axi_in_45_BREADY),
    .m_axi_BRESP(m_axi_in_45_BRESP),
    .m_axi_BVALID(m_axi_in_45_BVALID),
    .m_axi_RDATA(m_axi_in_45_RDATA),
    .m_axi_RID(m_axi_in_45_RID),
    .m_axi_RLAST(m_axi_in_45_RLAST),
    .m_axi_RREADY(m_axi_in_45_RREADY),
    .m_axi_RRESP(m_axi_in_45_RRESP),
    .m_axi_RVALID(m_axi_in_45_RVALID),
    .m_axi_WDATA(m_axi_in_45_WDATA),
    .m_axi_WLAST(m_axi_in_45_WLAST),
    .m_axi_WREADY(m_axi_in_45_WREADY),
    .m_axi_WSTRB(m_axi_in_45_WSTRB),
    .m_axi_WVALID(m_axi_in_45_WVALID),
    .read_addr_din(in_45_read_addr__din),
    .read_addr_full_n(in_45_read_addr__full_n),
    .read_addr_write(in_45_read_addr__write),
    .read_data_dout(in_45_read_data__dout),
    .read_data_empty_n(in_45_read_data__empty_n),
    .read_data_read(in_45_read_data__read),
    .write_addr_din(in_45_write_addr__din),
    .write_addr_full_n(in_45_write_addr__full_n),
    .write_addr_write(in_45_write_addr__write),
    .write_data_din(in_45_write_data__din),
    .write_data_full_n(in_45_write_data__full_n),
    .write_data_write(in_45_write_data__write),
    .write_resp_dout(in_45_write_resp__dout),
    .write_resp_empty_n(in_45_write_resp__empty_n),
    .write_resp_read(in_45_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_46__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_46_ARADDR),
    .m_axi_ARBURST(m_axi_in_46_ARBURST),
    .m_axi_ARCACHE(m_axi_in_46_ARCACHE),
    .m_axi_ARID(m_axi_in_46_ARID),
    .m_axi_ARLEN(m_axi_in_46_ARLEN),
    .m_axi_ARLOCK(m_axi_in_46_ARLOCK),
    .m_axi_ARPROT(m_axi_in_46_ARPROT),
    .m_axi_ARQOS(m_axi_in_46_ARQOS),
    .m_axi_ARREADY(m_axi_in_46_ARREADY),
    .m_axi_ARSIZE(m_axi_in_46_ARSIZE),
    .m_axi_ARVALID(m_axi_in_46_ARVALID),
    .m_axi_AWADDR(m_axi_in_46_AWADDR),
    .m_axi_AWBURST(m_axi_in_46_AWBURST),
    .m_axi_AWCACHE(m_axi_in_46_AWCACHE),
    .m_axi_AWID(m_axi_in_46_AWID),
    .m_axi_AWLEN(m_axi_in_46_AWLEN),
    .m_axi_AWLOCK(m_axi_in_46_AWLOCK),
    .m_axi_AWPROT(m_axi_in_46_AWPROT),
    .m_axi_AWQOS(m_axi_in_46_AWQOS),
    .m_axi_AWREADY(m_axi_in_46_AWREADY),
    .m_axi_AWSIZE(m_axi_in_46_AWSIZE),
    .m_axi_AWVALID(m_axi_in_46_AWVALID),
    .m_axi_BID(m_axi_in_46_BID),
    .m_axi_BREADY(m_axi_in_46_BREADY),
    .m_axi_BRESP(m_axi_in_46_BRESP),
    .m_axi_BVALID(m_axi_in_46_BVALID),
    .m_axi_RDATA(m_axi_in_46_RDATA),
    .m_axi_RID(m_axi_in_46_RID),
    .m_axi_RLAST(m_axi_in_46_RLAST),
    .m_axi_RREADY(m_axi_in_46_RREADY),
    .m_axi_RRESP(m_axi_in_46_RRESP),
    .m_axi_RVALID(m_axi_in_46_RVALID),
    .m_axi_WDATA(m_axi_in_46_WDATA),
    .m_axi_WLAST(m_axi_in_46_WLAST),
    .m_axi_WREADY(m_axi_in_46_WREADY),
    .m_axi_WSTRB(m_axi_in_46_WSTRB),
    .m_axi_WVALID(m_axi_in_46_WVALID),
    .read_addr_din(in_46_read_addr__din),
    .read_addr_full_n(in_46_read_addr__full_n),
    .read_addr_write(in_46_read_addr__write),
    .read_data_dout(in_46_read_data__dout),
    .read_data_empty_n(in_46_read_data__empty_n),
    .read_data_read(in_46_read_data__read),
    .write_addr_din(in_46_write_addr__din),
    .write_addr_full_n(in_46_write_addr__full_n),
    .write_addr_write(in_46_write_addr__write),
    .write_data_din(in_46_write_data__din),
    .write_data_full_n(in_46_write_data__full_n),
    .write_data_write(in_46_write_data__write),
    .write_resp_dout(in_46_write_resp__dout),
    .write_resp_empty_n(in_46_write_resp__empty_n),
    .write_resp_read(in_46_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_47__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_47_ARADDR),
    .m_axi_ARBURST(m_axi_in_47_ARBURST),
    .m_axi_ARCACHE(m_axi_in_47_ARCACHE),
    .m_axi_ARID(m_axi_in_47_ARID),
    .m_axi_ARLEN(m_axi_in_47_ARLEN),
    .m_axi_ARLOCK(m_axi_in_47_ARLOCK),
    .m_axi_ARPROT(m_axi_in_47_ARPROT),
    .m_axi_ARQOS(m_axi_in_47_ARQOS),
    .m_axi_ARREADY(m_axi_in_47_ARREADY),
    .m_axi_ARSIZE(m_axi_in_47_ARSIZE),
    .m_axi_ARVALID(m_axi_in_47_ARVALID),
    .m_axi_AWADDR(m_axi_in_47_AWADDR),
    .m_axi_AWBURST(m_axi_in_47_AWBURST),
    .m_axi_AWCACHE(m_axi_in_47_AWCACHE),
    .m_axi_AWID(m_axi_in_47_AWID),
    .m_axi_AWLEN(m_axi_in_47_AWLEN),
    .m_axi_AWLOCK(m_axi_in_47_AWLOCK),
    .m_axi_AWPROT(m_axi_in_47_AWPROT),
    .m_axi_AWQOS(m_axi_in_47_AWQOS),
    .m_axi_AWREADY(m_axi_in_47_AWREADY),
    .m_axi_AWSIZE(m_axi_in_47_AWSIZE),
    .m_axi_AWVALID(m_axi_in_47_AWVALID),
    .m_axi_BID(m_axi_in_47_BID),
    .m_axi_BREADY(m_axi_in_47_BREADY),
    .m_axi_BRESP(m_axi_in_47_BRESP),
    .m_axi_BVALID(m_axi_in_47_BVALID),
    .m_axi_RDATA(m_axi_in_47_RDATA),
    .m_axi_RID(m_axi_in_47_RID),
    .m_axi_RLAST(m_axi_in_47_RLAST),
    .m_axi_RREADY(m_axi_in_47_RREADY),
    .m_axi_RRESP(m_axi_in_47_RRESP),
    .m_axi_RVALID(m_axi_in_47_RVALID),
    .m_axi_WDATA(m_axi_in_47_WDATA),
    .m_axi_WLAST(m_axi_in_47_WLAST),
    .m_axi_WREADY(m_axi_in_47_WREADY),
    .m_axi_WSTRB(m_axi_in_47_WSTRB),
    .m_axi_WVALID(m_axi_in_47_WVALID),
    .read_addr_din(in_47_read_addr__din),
    .read_addr_full_n(in_47_read_addr__full_n),
    .read_addr_write(in_47_read_addr__write),
    .read_data_dout(in_47_read_data__dout),
    .read_data_empty_n(in_47_read_data__empty_n),
    .read_data_read(in_47_read_data__read),
    .write_addr_din(in_47_write_addr__din),
    .write_addr_full_n(in_47_write_addr__full_n),
    .write_addr_write(in_47_write_addr__write),
    .write_data_din(in_47_write_data__din),
    .write_data_full_n(in_47_write_data__full_n),
    .write_data_write(in_47_write_data__write),
    .write_resp_dout(in_47_write_resp__dout),
    .write_resp_empty_n(in_47_write_resp__empty_n),
    .write_resp_read(in_47_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_48__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_48_ARADDR),
    .m_axi_ARBURST(m_axi_in_48_ARBURST),
    .m_axi_ARCACHE(m_axi_in_48_ARCACHE),
    .m_axi_ARID(m_axi_in_48_ARID),
    .m_axi_ARLEN(m_axi_in_48_ARLEN),
    .m_axi_ARLOCK(m_axi_in_48_ARLOCK),
    .m_axi_ARPROT(m_axi_in_48_ARPROT),
    .m_axi_ARQOS(m_axi_in_48_ARQOS),
    .m_axi_ARREADY(m_axi_in_48_ARREADY),
    .m_axi_ARSIZE(m_axi_in_48_ARSIZE),
    .m_axi_ARVALID(m_axi_in_48_ARVALID),
    .m_axi_AWADDR(m_axi_in_48_AWADDR),
    .m_axi_AWBURST(m_axi_in_48_AWBURST),
    .m_axi_AWCACHE(m_axi_in_48_AWCACHE),
    .m_axi_AWID(m_axi_in_48_AWID),
    .m_axi_AWLEN(m_axi_in_48_AWLEN),
    .m_axi_AWLOCK(m_axi_in_48_AWLOCK),
    .m_axi_AWPROT(m_axi_in_48_AWPROT),
    .m_axi_AWQOS(m_axi_in_48_AWQOS),
    .m_axi_AWREADY(m_axi_in_48_AWREADY),
    .m_axi_AWSIZE(m_axi_in_48_AWSIZE),
    .m_axi_AWVALID(m_axi_in_48_AWVALID),
    .m_axi_BID(m_axi_in_48_BID),
    .m_axi_BREADY(m_axi_in_48_BREADY),
    .m_axi_BRESP(m_axi_in_48_BRESP),
    .m_axi_BVALID(m_axi_in_48_BVALID),
    .m_axi_RDATA(m_axi_in_48_RDATA),
    .m_axi_RID(m_axi_in_48_RID),
    .m_axi_RLAST(m_axi_in_48_RLAST),
    .m_axi_RREADY(m_axi_in_48_RREADY),
    .m_axi_RRESP(m_axi_in_48_RRESP),
    .m_axi_RVALID(m_axi_in_48_RVALID),
    .m_axi_WDATA(m_axi_in_48_WDATA),
    .m_axi_WLAST(m_axi_in_48_WLAST),
    .m_axi_WREADY(m_axi_in_48_WREADY),
    .m_axi_WSTRB(m_axi_in_48_WSTRB),
    .m_axi_WVALID(m_axi_in_48_WVALID),
    .read_addr_din(in_48_read_addr__din),
    .read_addr_full_n(in_48_read_addr__full_n),
    .read_addr_write(in_48_read_addr__write),
    .read_data_dout(in_48_read_data__dout),
    .read_data_empty_n(in_48_read_data__empty_n),
    .read_data_read(in_48_read_data__read),
    .write_addr_din(in_48_write_addr__din),
    .write_addr_full_n(in_48_write_addr__full_n),
    .write_addr_write(in_48_write_addr__write),
    .write_data_din(in_48_write_data__din),
    .write_data_full_n(in_48_write_data__full_n),
    .write_data_write(in_48_write_data__write),
    .write_resp_dout(in_48_write_resp__dout),
    .write_resp_empty_n(in_48_write_resp__empty_n),
    .write_resp_read(in_48_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_49__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_49_ARADDR),
    .m_axi_ARBURST(m_axi_in_49_ARBURST),
    .m_axi_ARCACHE(m_axi_in_49_ARCACHE),
    .m_axi_ARID(m_axi_in_49_ARID),
    .m_axi_ARLEN(m_axi_in_49_ARLEN),
    .m_axi_ARLOCK(m_axi_in_49_ARLOCK),
    .m_axi_ARPROT(m_axi_in_49_ARPROT),
    .m_axi_ARQOS(m_axi_in_49_ARQOS),
    .m_axi_ARREADY(m_axi_in_49_ARREADY),
    .m_axi_ARSIZE(m_axi_in_49_ARSIZE),
    .m_axi_ARVALID(m_axi_in_49_ARVALID),
    .m_axi_AWADDR(m_axi_in_49_AWADDR),
    .m_axi_AWBURST(m_axi_in_49_AWBURST),
    .m_axi_AWCACHE(m_axi_in_49_AWCACHE),
    .m_axi_AWID(m_axi_in_49_AWID),
    .m_axi_AWLEN(m_axi_in_49_AWLEN),
    .m_axi_AWLOCK(m_axi_in_49_AWLOCK),
    .m_axi_AWPROT(m_axi_in_49_AWPROT),
    .m_axi_AWQOS(m_axi_in_49_AWQOS),
    .m_axi_AWREADY(m_axi_in_49_AWREADY),
    .m_axi_AWSIZE(m_axi_in_49_AWSIZE),
    .m_axi_AWVALID(m_axi_in_49_AWVALID),
    .m_axi_BID(m_axi_in_49_BID),
    .m_axi_BREADY(m_axi_in_49_BREADY),
    .m_axi_BRESP(m_axi_in_49_BRESP),
    .m_axi_BVALID(m_axi_in_49_BVALID),
    .m_axi_RDATA(m_axi_in_49_RDATA),
    .m_axi_RID(m_axi_in_49_RID),
    .m_axi_RLAST(m_axi_in_49_RLAST),
    .m_axi_RREADY(m_axi_in_49_RREADY),
    .m_axi_RRESP(m_axi_in_49_RRESP),
    .m_axi_RVALID(m_axi_in_49_RVALID),
    .m_axi_WDATA(m_axi_in_49_WDATA),
    .m_axi_WLAST(m_axi_in_49_WLAST),
    .m_axi_WREADY(m_axi_in_49_WREADY),
    .m_axi_WSTRB(m_axi_in_49_WSTRB),
    .m_axi_WVALID(m_axi_in_49_WVALID),
    .read_addr_din(in_49_read_addr__din),
    .read_addr_full_n(in_49_read_addr__full_n),
    .read_addr_write(in_49_read_addr__write),
    .read_data_dout(in_49_read_data__dout),
    .read_data_empty_n(in_49_read_data__empty_n),
    .read_data_read(in_49_read_data__read),
    .write_addr_din(in_49_write_addr__din),
    .write_addr_full_n(in_49_write_addr__full_n),
    .write_addr_write(in_49_write_addr__write),
    .write_data_din(in_49_write_data__din),
    .write_data_full_n(in_49_write_data__full_n),
    .write_data_write(in_49_write_data__write),
    .write_resp_dout(in_49_write_resp__dout),
    .write_resp_empty_n(in_49_write_resp__empty_n),
    .write_resp_read(in_49_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_5_ARADDR),
    .m_axi_ARBURST(m_axi_in_5_ARBURST),
    .m_axi_ARCACHE(m_axi_in_5_ARCACHE),
    .m_axi_ARID(m_axi_in_5_ARID),
    .m_axi_ARLEN(m_axi_in_5_ARLEN),
    .m_axi_ARLOCK(m_axi_in_5_ARLOCK),
    .m_axi_ARPROT(m_axi_in_5_ARPROT),
    .m_axi_ARQOS(m_axi_in_5_ARQOS),
    .m_axi_ARREADY(m_axi_in_5_ARREADY),
    .m_axi_ARSIZE(m_axi_in_5_ARSIZE),
    .m_axi_ARVALID(m_axi_in_5_ARVALID),
    .m_axi_AWADDR(m_axi_in_5_AWADDR),
    .m_axi_AWBURST(m_axi_in_5_AWBURST),
    .m_axi_AWCACHE(m_axi_in_5_AWCACHE),
    .m_axi_AWID(m_axi_in_5_AWID),
    .m_axi_AWLEN(m_axi_in_5_AWLEN),
    .m_axi_AWLOCK(m_axi_in_5_AWLOCK),
    .m_axi_AWPROT(m_axi_in_5_AWPROT),
    .m_axi_AWQOS(m_axi_in_5_AWQOS),
    .m_axi_AWREADY(m_axi_in_5_AWREADY),
    .m_axi_AWSIZE(m_axi_in_5_AWSIZE),
    .m_axi_AWVALID(m_axi_in_5_AWVALID),
    .m_axi_BID(m_axi_in_5_BID),
    .m_axi_BREADY(m_axi_in_5_BREADY),
    .m_axi_BRESP(m_axi_in_5_BRESP),
    .m_axi_BVALID(m_axi_in_5_BVALID),
    .m_axi_RDATA(m_axi_in_5_RDATA),
    .m_axi_RID(m_axi_in_5_RID),
    .m_axi_RLAST(m_axi_in_5_RLAST),
    .m_axi_RREADY(m_axi_in_5_RREADY),
    .m_axi_RRESP(m_axi_in_5_RRESP),
    .m_axi_RVALID(m_axi_in_5_RVALID),
    .m_axi_WDATA(m_axi_in_5_WDATA),
    .m_axi_WLAST(m_axi_in_5_WLAST),
    .m_axi_WREADY(m_axi_in_5_WREADY),
    .m_axi_WSTRB(m_axi_in_5_WSTRB),
    .m_axi_WVALID(m_axi_in_5_WVALID),
    .read_addr_din(in_5_read_addr__din),
    .read_addr_full_n(in_5_read_addr__full_n),
    .read_addr_write(in_5_read_addr__write),
    .read_data_dout(in_5_read_data__dout),
    .read_data_empty_n(in_5_read_data__empty_n),
    .read_data_read(in_5_read_data__read),
    .write_addr_din(in_5_write_addr__din),
    .write_addr_full_n(in_5_write_addr__full_n),
    .write_addr_write(in_5_write_addr__write),
    .write_data_din(in_5_write_data__din),
    .write_data_full_n(in_5_write_data__full_n),
    .write_data_write(in_5_write_data__write),
    .write_resp_dout(in_5_write_resp__dout),
    .write_resp_empty_n(in_5_write_resp__empty_n),
    .write_resp_read(in_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_50__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_50_ARADDR),
    .m_axi_ARBURST(m_axi_in_50_ARBURST),
    .m_axi_ARCACHE(m_axi_in_50_ARCACHE),
    .m_axi_ARID(m_axi_in_50_ARID),
    .m_axi_ARLEN(m_axi_in_50_ARLEN),
    .m_axi_ARLOCK(m_axi_in_50_ARLOCK),
    .m_axi_ARPROT(m_axi_in_50_ARPROT),
    .m_axi_ARQOS(m_axi_in_50_ARQOS),
    .m_axi_ARREADY(m_axi_in_50_ARREADY),
    .m_axi_ARSIZE(m_axi_in_50_ARSIZE),
    .m_axi_ARVALID(m_axi_in_50_ARVALID),
    .m_axi_AWADDR(m_axi_in_50_AWADDR),
    .m_axi_AWBURST(m_axi_in_50_AWBURST),
    .m_axi_AWCACHE(m_axi_in_50_AWCACHE),
    .m_axi_AWID(m_axi_in_50_AWID),
    .m_axi_AWLEN(m_axi_in_50_AWLEN),
    .m_axi_AWLOCK(m_axi_in_50_AWLOCK),
    .m_axi_AWPROT(m_axi_in_50_AWPROT),
    .m_axi_AWQOS(m_axi_in_50_AWQOS),
    .m_axi_AWREADY(m_axi_in_50_AWREADY),
    .m_axi_AWSIZE(m_axi_in_50_AWSIZE),
    .m_axi_AWVALID(m_axi_in_50_AWVALID),
    .m_axi_BID(m_axi_in_50_BID),
    .m_axi_BREADY(m_axi_in_50_BREADY),
    .m_axi_BRESP(m_axi_in_50_BRESP),
    .m_axi_BVALID(m_axi_in_50_BVALID),
    .m_axi_RDATA(m_axi_in_50_RDATA),
    .m_axi_RID(m_axi_in_50_RID),
    .m_axi_RLAST(m_axi_in_50_RLAST),
    .m_axi_RREADY(m_axi_in_50_RREADY),
    .m_axi_RRESP(m_axi_in_50_RRESP),
    .m_axi_RVALID(m_axi_in_50_RVALID),
    .m_axi_WDATA(m_axi_in_50_WDATA),
    .m_axi_WLAST(m_axi_in_50_WLAST),
    .m_axi_WREADY(m_axi_in_50_WREADY),
    .m_axi_WSTRB(m_axi_in_50_WSTRB),
    .m_axi_WVALID(m_axi_in_50_WVALID),
    .read_addr_din(in_50_read_addr__din),
    .read_addr_full_n(in_50_read_addr__full_n),
    .read_addr_write(in_50_read_addr__write),
    .read_data_dout(in_50_read_data__dout),
    .read_data_empty_n(in_50_read_data__empty_n),
    .read_data_read(in_50_read_data__read),
    .write_addr_din(in_50_write_addr__din),
    .write_addr_full_n(in_50_write_addr__full_n),
    .write_addr_write(in_50_write_addr__write),
    .write_data_din(in_50_write_data__din),
    .write_data_full_n(in_50_write_data__full_n),
    .write_data_write(in_50_write_data__write),
    .write_resp_dout(in_50_write_resp__dout),
    .write_resp_empty_n(in_50_write_resp__empty_n),
    .write_resp_read(in_50_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_51__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_51_ARADDR),
    .m_axi_ARBURST(m_axi_in_51_ARBURST),
    .m_axi_ARCACHE(m_axi_in_51_ARCACHE),
    .m_axi_ARID(m_axi_in_51_ARID),
    .m_axi_ARLEN(m_axi_in_51_ARLEN),
    .m_axi_ARLOCK(m_axi_in_51_ARLOCK),
    .m_axi_ARPROT(m_axi_in_51_ARPROT),
    .m_axi_ARQOS(m_axi_in_51_ARQOS),
    .m_axi_ARREADY(m_axi_in_51_ARREADY),
    .m_axi_ARSIZE(m_axi_in_51_ARSIZE),
    .m_axi_ARVALID(m_axi_in_51_ARVALID),
    .m_axi_AWADDR(m_axi_in_51_AWADDR),
    .m_axi_AWBURST(m_axi_in_51_AWBURST),
    .m_axi_AWCACHE(m_axi_in_51_AWCACHE),
    .m_axi_AWID(m_axi_in_51_AWID),
    .m_axi_AWLEN(m_axi_in_51_AWLEN),
    .m_axi_AWLOCK(m_axi_in_51_AWLOCK),
    .m_axi_AWPROT(m_axi_in_51_AWPROT),
    .m_axi_AWQOS(m_axi_in_51_AWQOS),
    .m_axi_AWREADY(m_axi_in_51_AWREADY),
    .m_axi_AWSIZE(m_axi_in_51_AWSIZE),
    .m_axi_AWVALID(m_axi_in_51_AWVALID),
    .m_axi_BID(m_axi_in_51_BID),
    .m_axi_BREADY(m_axi_in_51_BREADY),
    .m_axi_BRESP(m_axi_in_51_BRESP),
    .m_axi_BVALID(m_axi_in_51_BVALID),
    .m_axi_RDATA(m_axi_in_51_RDATA),
    .m_axi_RID(m_axi_in_51_RID),
    .m_axi_RLAST(m_axi_in_51_RLAST),
    .m_axi_RREADY(m_axi_in_51_RREADY),
    .m_axi_RRESP(m_axi_in_51_RRESP),
    .m_axi_RVALID(m_axi_in_51_RVALID),
    .m_axi_WDATA(m_axi_in_51_WDATA),
    .m_axi_WLAST(m_axi_in_51_WLAST),
    .m_axi_WREADY(m_axi_in_51_WREADY),
    .m_axi_WSTRB(m_axi_in_51_WSTRB),
    .m_axi_WVALID(m_axi_in_51_WVALID),
    .read_addr_din(in_51_read_addr__din),
    .read_addr_full_n(in_51_read_addr__full_n),
    .read_addr_write(in_51_read_addr__write),
    .read_data_dout(in_51_read_data__dout),
    .read_data_empty_n(in_51_read_data__empty_n),
    .read_data_read(in_51_read_data__read),
    .write_addr_din(in_51_write_addr__din),
    .write_addr_full_n(in_51_write_addr__full_n),
    .write_addr_write(in_51_write_addr__write),
    .write_data_din(in_51_write_data__din),
    .write_data_full_n(in_51_write_data__full_n),
    .write_data_write(in_51_write_data__write),
    .write_resp_dout(in_51_write_resp__dout),
    .write_resp_empty_n(in_51_write_resp__empty_n),
    .write_resp_read(in_51_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_52__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_52_ARADDR),
    .m_axi_ARBURST(m_axi_in_52_ARBURST),
    .m_axi_ARCACHE(m_axi_in_52_ARCACHE),
    .m_axi_ARID(m_axi_in_52_ARID),
    .m_axi_ARLEN(m_axi_in_52_ARLEN),
    .m_axi_ARLOCK(m_axi_in_52_ARLOCK),
    .m_axi_ARPROT(m_axi_in_52_ARPROT),
    .m_axi_ARQOS(m_axi_in_52_ARQOS),
    .m_axi_ARREADY(m_axi_in_52_ARREADY),
    .m_axi_ARSIZE(m_axi_in_52_ARSIZE),
    .m_axi_ARVALID(m_axi_in_52_ARVALID),
    .m_axi_AWADDR(m_axi_in_52_AWADDR),
    .m_axi_AWBURST(m_axi_in_52_AWBURST),
    .m_axi_AWCACHE(m_axi_in_52_AWCACHE),
    .m_axi_AWID(m_axi_in_52_AWID),
    .m_axi_AWLEN(m_axi_in_52_AWLEN),
    .m_axi_AWLOCK(m_axi_in_52_AWLOCK),
    .m_axi_AWPROT(m_axi_in_52_AWPROT),
    .m_axi_AWQOS(m_axi_in_52_AWQOS),
    .m_axi_AWREADY(m_axi_in_52_AWREADY),
    .m_axi_AWSIZE(m_axi_in_52_AWSIZE),
    .m_axi_AWVALID(m_axi_in_52_AWVALID),
    .m_axi_BID(m_axi_in_52_BID),
    .m_axi_BREADY(m_axi_in_52_BREADY),
    .m_axi_BRESP(m_axi_in_52_BRESP),
    .m_axi_BVALID(m_axi_in_52_BVALID),
    .m_axi_RDATA(m_axi_in_52_RDATA),
    .m_axi_RID(m_axi_in_52_RID),
    .m_axi_RLAST(m_axi_in_52_RLAST),
    .m_axi_RREADY(m_axi_in_52_RREADY),
    .m_axi_RRESP(m_axi_in_52_RRESP),
    .m_axi_RVALID(m_axi_in_52_RVALID),
    .m_axi_WDATA(m_axi_in_52_WDATA),
    .m_axi_WLAST(m_axi_in_52_WLAST),
    .m_axi_WREADY(m_axi_in_52_WREADY),
    .m_axi_WSTRB(m_axi_in_52_WSTRB),
    .m_axi_WVALID(m_axi_in_52_WVALID),
    .read_addr_din(in_52_read_addr__din),
    .read_addr_full_n(in_52_read_addr__full_n),
    .read_addr_write(in_52_read_addr__write),
    .read_data_dout(in_52_read_data__dout),
    .read_data_empty_n(in_52_read_data__empty_n),
    .read_data_read(in_52_read_data__read),
    .write_addr_din(in_52_write_addr__din),
    .write_addr_full_n(in_52_write_addr__full_n),
    .write_addr_write(in_52_write_addr__write),
    .write_data_din(in_52_write_data__din),
    .write_data_full_n(in_52_write_data__full_n),
    .write_data_write(in_52_write_data__write),
    .write_resp_dout(in_52_write_resp__dout),
    .write_resp_empty_n(in_52_write_resp__empty_n),
    .write_resp_read(in_52_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_53__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_53_ARADDR),
    .m_axi_ARBURST(m_axi_in_53_ARBURST),
    .m_axi_ARCACHE(m_axi_in_53_ARCACHE),
    .m_axi_ARID(m_axi_in_53_ARID),
    .m_axi_ARLEN(m_axi_in_53_ARLEN),
    .m_axi_ARLOCK(m_axi_in_53_ARLOCK),
    .m_axi_ARPROT(m_axi_in_53_ARPROT),
    .m_axi_ARQOS(m_axi_in_53_ARQOS),
    .m_axi_ARREADY(m_axi_in_53_ARREADY),
    .m_axi_ARSIZE(m_axi_in_53_ARSIZE),
    .m_axi_ARVALID(m_axi_in_53_ARVALID),
    .m_axi_AWADDR(m_axi_in_53_AWADDR),
    .m_axi_AWBURST(m_axi_in_53_AWBURST),
    .m_axi_AWCACHE(m_axi_in_53_AWCACHE),
    .m_axi_AWID(m_axi_in_53_AWID),
    .m_axi_AWLEN(m_axi_in_53_AWLEN),
    .m_axi_AWLOCK(m_axi_in_53_AWLOCK),
    .m_axi_AWPROT(m_axi_in_53_AWPROT),
    .m_axi_AWQOS(m_axi_in_53_AWQOS),
    .m_axi_AWREADY(m_axi_in_53_AWREADY),
    .m_axi_AWSIZE(m_axi_in_53_AWSIZE),
    .m_axi_AWVALID(m_axi_in_53_AWVALID),
    .m_axi_BID(m_axi_in_53_BID),
    .m_axi_BREADY(m_axi_in_53_BREADY),
    .m_axi_BRESP(m_axi_in_53_BRESP),
    .m_axi_BVALID(m_axi_in_53_BVALID),
    .m_axi_RDATA(m_axi_in_53_RDATA),
    .m_axi_RID(m_axi_in_53_RID),
    .m_axi_RLAST(m_axi_in_53_RLAST),
    .m_axi_RREADY(m_axi_in_53_RREADY),
    .m_axi_RRESP(m_axi_in_53_RRESP),
    .m_axi_RVALID(m_axi_in_53_RVALID),
    .m_axi_WDATA(m_axi_in_53_WDATA),
    .m_axi_WLAST(m_axi_in_53_WLAST),
    .m_axi_WREADY(m_axi_in_53_WREADY),
    .m_axi_WSTRB(m_axi_in_53_WSTRB),
    .m_axi_WVALID(m_axi_in_53_WVALID),
    .read_addr_din(in_53_read_addr__din),
    .read_addr_full_n(in_53_read_addr__full_n),
    .read_addr_write(in_53_read_addr__write),
    .read_data_dout(in_53_read_data__dout),
    .read_data_empty_n(in_53_read_data__empty_n),
    .read_data_read(in_53_read_data__read),
    .write_addr_din(in_53_write_addr__din),
    .write_addr_full_n(in_53_write_addr__full_n),
    .write_addr_write(in_53_write_addr__write),
    .write_data_din(in_53_write_data__din),
    .write_data_full_n(in_53_write_data__full_n),
    .write_data_write(in_53_write_data__write),
    .write_resp_dout(in_53_write_resp__dout),
    .write_resp_empty_n(in_53_write_resp__empty_n),
    .write_resp_read(in_53_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_6_ARADDR),
    .m_axi_ARBURST(m_axi_in_6_ARBURST),
    .m_axi_ARCACHE(m_axi_in_6_ARCACHE),
    .m_axi_ARID(m_axi_in_6_ARID),
    .m_axi_ARLEN(m_axi_in_6_ARLEN),
    .m_axi_ARLOCK(m_axi_in_6_ARLOCK),
    .m_axi_ARPROT(m_axi_in_6_ARPROT),
    .m_axi_ARQOS(m_axi_in_6_ARQOS),
    .m_axi_ARREADY(m_axi_in_6_ARREADY),
    .m_axi_ARSIZE(m_axi_in_6_ARSIZE),
    .m_axi_ARVALID(m_axi_in_6_ARVALID),
    .m_axi_AWADDR(m_axi_in_6_AWADDR),
    .m_axi_AWBURST(m_axi_in_6_AWBURST),
    .m_axi_AWCACHE(m_axi_in_6_AWCACHE),
    .m_axi_AWID(m_axi_in_6_AWID),
    .m_axi_AWLEN(m_axi_in_6_AWLEN),
    .m_axi_AWLOCK(m_axi_in_6_AWLOCK),
    .m_axi_AWPROT(m_axi_in_6_AWPROT),
    .m_axi_AWQOS(m_axi_in_6_AWQOS),
    .m_axi_AWREADY(m_axi_in_6_AWREADY),
    .m_axi_AWSIZE(m_axi_in_6_AWSIZE),
    .m_axi_AWVALID(m_axi_in_6_AWVALID),
    .m_axi_BID(m_axi_in_6_BID),
    .m_axi_BREADY(m_axi_in_6_BREADY),
    .m_axi_BRESP(m_axi_in_6_BRESP),
    .m_axi_BVALID(m_axi_in_6_BVALID),
    .m_axi_RDATA(m_axi_in_6_RDATA),
    .m_axi_RID(m_axi_in_6_RID),
    .m_axi_RLAST(m_axi_in_6_RLAST),
    .m_axi_RREADY(m_axi_in_6_RREADY),
    .m_axi_RRESP(m_axi_in_6_RRESP),
    .m_axi_RVALID(m_axi_in_6_RVALID),
    .m_axi_WDATA(m_axi_in_6_WDATA),
    .m_axi_WLAST(m_axi_in_6_WLAST),
    .m_axi_WREADY(m_axi_in_6_WREADY),
    .m_axi_WSTRB(m_axi_in_6_WSTRB),
    .m_axi_WVALID(m_axi_in_6_WVALID),
    .read_addr_din(in_6_read_addr__din),
    .read_addr_full_n(in_6_read_addr__full_n),
    .read_addr_write(in_6_read_addr__write),
    .read_data_dout(in_6_read_data__dout),
    .read_data_empty_n(in_6_read_data__empty_n),
    .read_data_read(in_6_read_data__read),
    .write_addr_din(in_6_write_addr__din),
    .write_addr_full_n(in_6_write_addr__full_n),
    .write_addr_write(in_6_write_addr__write),
    .write_data_din(in_6_write_data__din),
    .write_data_full_n(in_6_write_data__full_n),
    .write_data_write(in_6_write_data__write),
    .write_resp_dout(in_6_write_resp__dout),
    .write_resp_empty_n(in_6_write_resp__empty_n),
    .write_resp_read(in_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_7_ARADDR),
    .m_axi_ARBURST(m_axi_in_7_ARBURST),
    .m_axi_ARCACHE(m_axi_in_7_ARCACHE),
    .m_axi_ARID(m_axi_in_7_ARID),
    .m_axi_ARLEN(m_axi_in_7_ARLEN),
    .m_axi_ARLOCK(m_axi_in_7_ARLOCK),
    .m_axi_ARPROT(m_axi_in_7_ARPROT),
    .m_axi_ARQOS(m_axi_in_7_ARQOS),
    .m_axi_ARREADY(m_axi_in_7_ARREADY),
    .m_axi_ARSIZE(m_axi_in_7_ARSIZE),
    .m_axi_ARVALID(m_axi_in_7_ARVALID),
    .m_axi_AWADDR(m_axi_in_7_AWADDR),
    .m_axi_AWBURST(m_axi_in_7_AWBURST),
    .m_axi_AWCACHE(m_axi_in_7_AWCACHE),
    .m_axi_AWID(m_axi_in_7_AWID),
    .m_axi_AWLEN(m_axi_in_7_AWLEN),
    .m_axi_AWLOCK(m_axi_in_7_AWLOCK),
    .m_axi_AWPROT(m_axi_in_7_AWPROT),
    .m_axi_AWQOS(m_axi_in_7_AWQOS),
    .m_axi_AWREADY(m_axi_in_7_AWREADY),
    .m_axi_AWSIZE(m_axi_in_7_AWSIZE),
    .m_axi_AWVALID(m_axi_in_7_AWVALID),
    .m_axi_BID(m_axi_in_7_BID),
    .m_axi_BREADY(m_axi_in_7_BREADY),
    .m_axi_BRESP(m_axi_in_7_BRESP),
    .m_axi_BVALID(m_axi_in_7_BVALID),
    .m_axi_RDATA(m_axi_in_7_RDATA),
    .m_axi_RID(m_axi_in_7_RID),
    .m_axi_RLAST(m_axi_in_7_RLAST),
    .m_axi_RREADY(m_axi_in_7_RREADY),
    .m_axi_RRESP(m_axi_in_7_RRESP),
    .m_axi_RVALID(m_axi_in_7_RVALID),
    .m_axi_WDATA(m_axi_in_7_WDATA),
    .m_axi_WLAST(m_axi_in_7_WLAST),
    .m_axi_WREADY(m_axi_in_7_WREADY),
    .m_axi_WSTRB(m_axi_in_7_WSTRB),
    .m_axi_WVALID(m_axi_in_7_WVALID),
    .read_addr_din(in_7_read_addr__din),
    .read_addr_full_n(in_7_read_addr__full_n),
    .read_addr_write(in_7_read_addr__write),
    .read_data_dout(in_7_read_data__dout),
    .read_data_empty_n(in_7_read_data__empty_n),
    .read_data_read(in_7_read_data__read),
    .write_addr_din(in_7_write_addr__din),
    .write_addr_full_n(in_7_write_addr__full_n),
    .write_addr_write(in_7_write_addr__write),
    .write_data_din(in_7_write_data__din),
    .write_data_full_n(in_7_write_data__full_n),
    .write_data_write(in_7_write_data__write),
    .write_resp_dout(in_7_write_resp__dout),
    .write_resp_empty_n(in_7_write_resp__empty_n),
    .write_resp_read(in_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_8__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_8_ARADDR),
    .m_axi_ARBURST(m_axi_in_8_ARBURST),
    .m_axi_ARCACHE(m_axi_in_8_ARCACHE),
    .m_axi_ARID(m_axi_in_8_ARID),
    .m_axi_ARLEN(m_axi_in_8_ARLEN),
    .m_axi_ARLOCK(m_axi_in_8_ARLOCK),
    .m_axi_ARPROT(m_axi_in_8_ARPROT),
    .m_axi_ARQOS(m_axi_in_8_ARQOS),
    .m_axi_ARREADY(m_axi_in_8_ARREADY),
    .m_axi_ARSIZE(m_axi_in_8_ARSIZE),
    .m_axi_ARVALID(m_axi_in_8_ARVALID),
    .m_axi_AWADDR(m_axi_in_8_AWADDR),
    .m_axi_AWBURST(m_axi_in_8_AWBURST),
    .m_axi_AWCACHE(m_axi_in_8_AWCACHE),
    .m_axi_AWID(m_axi_in_8_AWID),
    .m_axi_AWLEN(m_axi_in_8_AWLEN),
    .m_axi_AWLOCK(m_axi_in_8_AWLOCK),
    .m_axi_AWPROT(m_axi_in_8_AWPROT),
    .m_axi_AWQOS(m_axi_in_8_AWQOS),
    .m_axi_AWREADY(m_axi_in_8_AWREADY),
    .m_axi_AWSIZE(m_axi_in_8_AWSIZE),
    .m_axi_AWVALID(m_axi_in_8_AWVALID),
    .m_axi_BID(m_axi_in_8_BID),
    .m_axi_BREADY(m_axi_in_8_BREADY),
    .m_axi_BRESP(m_axi_in_8_BRESP),
    .m_axi_BVALID(m_axi_in_8_BVALID),
    .m_axi_RDATA(m_axi_in_8_RDATA),
    .m_axi_RID(m_axi_in_8_RID),
    .m_axi_RLAST(m_axi_in_8_RLAST),
    .m_axi_RREADY(m_axi_in_8_RREADY),
    .m_axi_RRESP(m_axi_in_8_RRESP),
    .m_axi_RVALID(m_axi_in_8_RVALID),
    .m_axi_WDATA(m_axi_in_8_WDATA),
    .m_axi_WLAST(m_axi_in_8_WLAST),
    .m_axi_WREADY(m_axi_in_8_WREADY),
    .m_axi_WSTRB(m_axi_in_8_WSTRB),
    .m_axi_WVALID(m_axi_in_8_WVALID),
    .read_addr_din(in_8_read_addr__din),
    .read_addr_full_n(in_8_read_addr__full_n),
    .read_addr_write(in_8_read_addr__write),
    .read_data_dout(in_8_read_data__dout),
    .read_data_empty_n(in_8_read_data__empty_n),
    .read_data_read(in_8_read_data__read),
    .write_addr_din(in_8_write_addr__din),
    .write_addr_full_n(in_8_write_addr__full_n),
    .write_addr_write(in_8_write_addr__write),
    .write_data_din(in_8_write_data__din),
    .write_data_full_n(in_8_write_data__full_n),
    .write_data_write(in_8_write_data__write),
    .write_resp_dout(in_8_write_resp__dout),
    .write_resp_empty_n(in_8_write_resp__empty_n),
    .write_resp_read(in_8_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_9__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_9_ARADDR),
    .m_axi_ARBURST(m_axi_in_9_ARBURST),
    .m_axi_ARCACHE(m_axi_in_9_ARCACHE),
    .m_axi_ARID(m_axi_in_9_ARID),
    .m_axi_ARLEN(m_axi_in_9_ARLEN),
    .m_axi_ARLOCK(m_axi_in_9_ARLOCK),
    .m_axi_ARPROT(m_axi_in_9_ARPROT),
    .m_axi_ARQOS(m_axi_in_9_ARQOS),
    .m_axi_ARREADY(m_axi_in_9_ARREADY),
    .m_axi_ARSIZE(m_axi_in_9_ARSIZE),
    .m_axi_ARVALID(m_axi_in_9_ARVALID),
    .m_axi_AWADDR(m_axi_in_9_AWADDR),
    .m_axi_AWBURST(m_axi_in_9_AWBURST),
    .m_axi_AWCACHE(m_axi_in_9_AWCACHE),
    .m_axi_AWID(m_axi_in_9_AWID),
    .m_axi_AWLEN(m_axi_in_9_AWLEN),
    .m_axi_AWLOCK(m_axi_in_9_AWLOCK),
    .m_axi_AWPROT(m_axi_in_9_AWPROT),
    .m_axi_AWQOS(m_axi_in_9_AWQOS),
    .m_axi_AWREADY(m_axi_in_9_AWREADY),
    .m_axi_AWSIZE(m_axi_in_9_AWSIZE),
    .m_axi_AWVALID(m_axi_in_9_AWVALID),
    .m_axi_BID(m_axi_in_9_BID),
    .m_axi_BREADY(m_axi_in_9_BREADY),
    .m_axi_BRESP(m_axi_in_9_BRESP),
    .m_axi_BVALID(m_axi_in_9_BVALID),
    .m_axi_RDATA(m_axi_in_9_RDATA),
    .m_axi_RID(m_axi_in_9_RID),
    .m_axi_RLAST(m_axi_in_9_RLAST),
    .m_axi_RREADY(m_axi_in_9_RREADY),
    .m_axi_RRESP(m_axi_in_9_RRESP),
    .m_axi_RVALID(m_axi_in_9_RVALID),
    .m_axi_WDATA(m_axi_in_9_WDATA),
    .m_axi_WLAST(m_axi_in_9_WLAST),
    .m_axi_WREADY(m_axi_in_9_WREADY),
    .m_axi_WSTRB(m_axi_in_9_WSTRB),
    .m_axi_WVALID(m_axi_in_9_WVALID),
    .read_addr_din(in_9_read_addr__din),
    .read_addr_full_n(in_9_read_addr__full_n),
    .read_addr_write(in_9_read_addr__write),
    .read_data_dout(in_9_read_data__dout),
    .read_data_empty_n(in_9_read_data__empty_n),
    .read_data_read(in_9_read_data__read),
    .write_addr_din(in_9_write_addr__din),
    .write_addr_full_n(in_9_write_addr__full_n),
    .write_addr_write(in_9_write_addr__write),
    .write_data_din(in_9_write_data__din),
    .write_data_full_n(in_9_write_data__full_n),
    .write_data_write(in_9_write_data__write),
    .write_resp_dout(in_9_write_resp__dout),
    .write_resp_empty_n(in_9_write_resp__empty_n),
    .write_resp_read(in_9_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) Knn_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .L4_out_dist(L4_out_dist),
    .L4_out_id(L4_out_id),
    .in_0(in_0),
    .in_1(in_1),
    .in_10(in_10),
    .in_11(in_11),
    .in_12(in_12),
    .in_13(in_13),
    .in_14(in_14),
    .in_15(in_15),
    .in_16(in_16),
    .in_17(in_17),
    .in_18(in_18),
    .in_19(in_19),
    .in_2(in_2),
    .in_20(in_20),
    .in_21(in_21),
    .in_22(in_22),
    .in_23(in_23),
    .in_24(in_24),
    .in_25(in_25),
    .in_26(in_26),
    .in_27(in_27),
    .in_28(in_28),
    .in_29(in_29),
    .in_3(in_3),
    .in_30(in_30),
    .in_31(in_31),
    .in_32(in_32),
    .in_33(in_33),
    .in_34(in_34),
    .in_35(in_35),
    .in_36(in_36),
    .in_37(in_37),
    .in_38(in_38),
    .in_39(in_39),
    .in_4(in_4),
    .in_40(in_40),
    .in_41(in_41),
    .in_42(in_42),
    .in_43(in_43),
    .in_44(in_44),
    .in_45(in_45),
    .in_46(in_46),
    .in_47(in_47),
    .in_48(in_48),
    .in_49(in_49),
    .in_5(in_5),
    .in_50(in_50),
    .in_51(in_51),
    .in_52(in_52),
    .in_53(in_53),
    .in_6(in_6),
    .in_7(in_7),
    .in_8(in_8),
    .in_9(in_9),
    .krnl_globalSort_L1_L2_0__ap_start(krnl_globalSort_L1_L2_0__ap_start),
    .krnl_globalSort_L1_L2_0__ap_ready(krnl_globalSort_L1_L2_0__ap_ready),
    .krnl_globalSort_L1_L2_0__ap_done(krnl_globalSort_L1_L2_0__ap_done),
    .krnl_globalSort_L1_L2_0__ap_idle(krnl_globalSort_L1_L2_0__ap_idle),
    .krnl_globalSort_L1_L2_1__ap_start(krnl_globalSort_L1_L2_1__ap_start),
    .krnl_globalSort_L1_L2_1__ap_ready(krnl_globalSort_L1_L2_1__ap_ready),
    .krnl_globalSort_L1_L2_1__ap_done(krnl_globalSort_L1_L2_1__ap_done),
    .krnl_globalSort_L1_L2_1__ap_idle(krnl_globalSort_L1_L2_1__ap_idle),
    .krnl_globalSort_L1_L2_2__ap_start(krnl_globalSort_L1_L2_2__ap_start),
    .krnl_globalSort_L1_L2_2__ap_ready(krnl_globalSort_L1_L2_2__ap_ready),
    .krnl_globalSort_L1_L2_2__ap_done(krnl_globalSort_L1_L2_2__ap_done),
    .krnl_globalSort_L1_L2_2__ap_idle(krnl_globalSort_L1_L2_2__ap_idle),
    .krnl_globalSort_L1_L2_3__ap_start(krnl_globalSort_L1_L2_3__ap_start),
    .krnl_globalSort_L1_L2_3__ap_ready(krnl_globalSort_L1_L2_3__ap_ready),
    .krnl_globalSort_L1_L2_3__ap_done(krnl_globalSort_L1_L2_3__ap_done),
    .krnl_globalSort_L1_L2_3__ap_idle(krnl_globalSort_L1_L2_3__ap_idle),
    .krnl_globalSort_L1_L2_4__ap_start(krnl_globalSort_L1_L2_4__ap_start),
    .krnl_globalSort_L1_L2_4__ap_ready(krnl_globalSort_L1_L2_4__ap_ready),
    .krnl_globalSort_L1_L2_4__ap_done(krnl_globalSort_L1_L2_4__ap_done),
    .krnl_globalSort_L1_L2_4__ap_idle(krnl_globalSort_L1_L2_4__ap_idle),
    .krnl_globalSort_L1_L2_5__ap_start(krnl_globalSort_L1_L2_5__ap_start),
    .krnl_globalSort_L1_L2_5__ap_ready(krnl_globalSort_L1_L2_5__ap_ready),
    .krnl_globalSort_L1_L2_5__ap_done(krnl_globalSort_L1_L2_5__ap_done),
    .krnl_globalSort_L1_L2_5__ap_idle(krnl_globalSort_L1_L2_5__ap_idle),
    .krnl_globalSort_L1_L2_6__ap_start(krnl_globalSort_L1_L2_6__ap_start),
    .krnl_globalSort_L1_L2_6__ap_ready(krnl_globalSort_L1_L2_6__ap_ready),
    .krnl_globalSort_L1_L2_6__ap_done(krnl_globalSort_L1_L2_6__ap_done),
    .krnl_globalSort_L1_L2_6__ap_idle(krnl_globalSort_L1_L2_6__ap_idle),
    .krnl_globalSort_L1_L2_7__ap_start(krnl_globalSort_L1_L2_7__ap_start),
    .krnl_globalSort_L1_L2_7__ap_ready(krnl_globalSort_L1_L2_7__ap_ready),
    .krnl_globalSort_L1_L2_7__ap_done(krnl_globalSort_L1_L2_7__ap_done),
    .krnl_globalSort_L1_L2_7__ap_idle(krnl_globalSort_L1_L2_7__ap_idle),
    .krnl_globalSort_L1_L2_8__ap_start(krnl_globalSort_L1_L2_8__ap_start),
    .krnl_globalSort_L1_L2_8__ap_ready(krnl_globalSort_L1_L2_8__ap_ready),
    .krnl_globalSort_L1_L2_8__ap_done(krnl_globalSort_L1_L2_8__ap_done),
    .krnl_globalSort_L1_L2_8__ap_idle(krnl_globalSort_L1_L2_8__ap_idle),
    .krnl_globalSort_L1_L2_9__ap_start(krnl_globalSort_L1_L2_9__ap_start),
    .krnl_globalSort_L1_L2_9__ap_ready(krnl_globalSort_L1_L2_9__ap_ready),
    .krnl_globalSort_L1_L2_9__ap_done(krnl_globalSort_L1_L2_9__ap_done),
    .krnl_globalSort_L1_L2_9__ap_idle(krnl_globalSort_L1_L2_9__ap_idle),
    .krnl_globalSort_L1_L2_10__ap_start(krnl_globalSort_L1_L2_10__ap_start),
    .krnl_globalSort_L1_L2_10__ap_ready(krnl_globalSort_L1_L2_10__ap_ready),
    .krnl_globalSort_L1_L2_10__ap_done(krnl_globalSort_L1_L2_10__ap_done),
    .krnl_globalSort_L1_L2_10__ap_idle(krnl_globalSort_L1_L2_10__ap_idle),
    .krnl_globalSort_L1_L2_11__ap_start(krnl_globalSort_L1_L2_11__ap_start),
    .krnl_globalSort_L1_L2_11__ap_ready(krnl_globalSort_L1_L2_11__ap_ready),
    .krnl_globalSort_L1_L2_11__ap_done(krnl_globalSort_L1_L2_11__ap_done),
    .krnl_globalSort_L1_L2_11__ap_idle(krnl_globalSort_L1_L2_11__ap_idle),
    .krnl_globalSort_L1_L2_12__ap_start(krnl_globalSort_L1_L2_12__ap_start),
    .krnl_globalSort_L1_L2_12__ap_ready(krnl_globalSort_L1_L2_12__ap_ready),
    .krnl_globalSort_L1_L2_12__ap_done(krnl_globalSort_L1_L2_12__ap_done),
    .krnl_globalSort_L1_L2_12__ap_idle(krnl_globalSort_L1_L2_12__ap_idle),
    .krnl_globalSort_L1_L2_13__ap_start(krnl_globalSort_L1_L2_13__ap_start),
    .krnl_globalSort_L1_L2_13__ap_ready(krnl_globalSort_L1_L2_13__ap_ready),
    .krnl_globalSort_L1_L2_13__ap_done(krnl_globalSort_L1_L2_13__ap_done),
    .krnl_globalSort_L1_L2_13__ap_idle(krnl_globalSort_L1_L2_13__ap_idle),
    .krnl_globalSort_L1_L2_14__ap_start(krnl_globalSort_L1_L2_14__ap_start),
    .krnl_globalSort_L1_L2_14__ap_ready(krnl_globalSort_L1_L2_14__ap_ready),
    .krnl_globalSort_L1_L2_14__ap_done(krnl_globalSort_L1_L2_14__ap_done),
    .krnl_globalSort_L1_L2_14__ap_idle(krnl_globalSort_L1_L2_14__ap_idle),
    .krnl_globalSort_L1_L2_15__ap_start(krnl_globalSort_L1_L2_15__ap_start),
    .krnl_globalSort_L1_L2_15__ap_ready(krnl_globalSort_L1_L2_15__ap_ready),
    .krnl_globalSort_L1_L2_15__ap_done(krnl_globalSort_L1_L2_15__ap_done),
    .krnl_globalSort_L1_L2_15__ap_idle(krnl_globalSort_L1_L2_15__ap_idle),
    .krnl_globalSort_L1_L2_16__ap_start(krnl_globalSort_L1_L2_16__ap_start),
    .krnl_globalSort_L1_L2_16__ap_ready(krnl_globalSort_L1_L2_16__ap_ready),
    .krnl_globalSort_L1_L2_16__ap_done(krnl_globalSort_L1_L2_16__ap_done),
    .krnl_globalSort_L1_L2_16__ap_idle(krnl_globalSort_L1_L2_16__ap_idle),
    .krnl_globalSort_L1_L2_17__ap_start(krnl_globalSort_L1_L2_17__ap_start),
    .krnl_globalSort_L1_L2_17__ap_ready(krnl_globalSort_L1_L2_17__ap_ready),
    .krnl_globalSort_L1_L2_17__ap_done(krnl_globalSort_L1_L2_17__ap_done),
    .krnl_globalSort_L1_L2_17__ap_idle(krnl_globalSort_L1_L2_17__ap_idle),
    .krnl_globalSort_L1_L2_18__ap_start(krnl_globalSort_L1_L2_18__ap_start),
    .krnl_globalSort_L1_L2_18__ap_ready(krnl_globalSort_L1_L2_18__ap_ready),
    .krnl_globalSort_L1_L2_18__ap_done(krnl_globalSort_L1_L2_18__ap_done),
    .krnl_globalSort_L1_L2_18__ap_idle(krnl_globalSort_L1_L2_18__ap_idle),
    .krnl_globalSort_L1_L2_19__ap_start(krnl_globalSort_L1_L2_19__ap_start),
    .krnl_globalSort_L1_L2_19__ap_ready(krnl_globalSort_L1_L2_19__ap_ready),
    .krnl_globalSort_L1_L2_19__ap_done(krnl_globalSort_L1_L2_19__ap_done),
    .krnl_globalSort_L1_L2_19__ap_idle(krnl_globalSort_L1_L2_19__ap_idle),
    .krnl_globalSort_L1_L2_20__ap_start(krnl_globalSort_L1_L2_20__ap_start),
    .krnl_globalSort_L1_L2_20__ap_ready(krnl_globalSort_L1_L2_20__ap_ready),
    .krnl_globalSort_L1_L2_20__ap_done(krnl_globalSort_L1_L2_20__ap_done),
    .krnl_globalSort_L1_L2_20__ap_idle(krnl_globalSort_L1_L2_20__ap_idle),
    .krnl_globalSort_L1_L2_21__ap_start(krnl_globalSort_L1_L2_21__ap_start),
    .krnl_globalSort_L1_L2_21__ap_ready(krnl_globalSort_L1_L2_21__ap_ready),
    .krnl_globalSort_L1_L2_21__ap_done(krnl_globalSort_L1_L2_21__ap_done),
    .krnl_globalSort_L1_L2_21__ap_idle(krnl_globalSort_L1_L2_21__ap_idle),
    .krnl_globalSort_L1_L2_22__ap_start(krnl_globalSort_L1_L2_22__ap_start),
    .krnl_globalSort_L1_L2_22__ap_ready(krnl_globalSort_L1_L2_22__ap_ready),
    .krnl_globalSort_L1_L2_22__ap_done(krnl_globalSort_L1_L2_22__ap_done),
    .krnl_globalSort_L1_L2_22__ap_idle(krnl_globalSort_L1_L2_22__ap_idle),
    .krnl_globalSort_L1_L2_23__ap_start(krnl_globalSort_L1_L2_23__ap_start),
    .krnl_globalSort_L1_L2_23__ap_ready(krnl_globalSort_L1_L2_23__ap_ready),
    .krnl_globalSort_L1_L2_23__ap_done(krnl_globalSort_L1_L2_23__ap_done),
    .krnl_globalSort_L1_L2_23__ap_idle(krnl_globalSort_L1_L2_23__ap_idle),
    .krnl_globalSort_L1_L2_24__ap_start(krnl_globalSort_L1_L2_24__ap_start),
    .krnl_globalSort_L1_L2_24__ap_ready(krnl_globalSort_L1_L2_24__ap_ready),
    .krnl_globalSort_L1_L2_24__ap_done(krnl_globalSort_L1_L2_24__ap_done),
    .krnl_globalSort_L1_L2_24__ap_idle(krnl_globalSort_L1_L2_24__ap_idle),
    .krnl_globalSort_L1_L2_25__ap_start(krnl_globalSort_L1_L2_25__ap_start),
    .krnl_globalSort_L1_L2_25__ap_ready(krnl_globalSort_L1_L2_25__ap_ready),
    .krnl_globalSort_L1_L2_25__ap_done(krnl_globalSort_L1_L2_25__ap_done),
    .krnl_globalSort_L1_L2_25__ap_idle(krnl_globalSort_L1_L2_25__ap_idle),
    .krnl_globalSort_L3_0___L4_out_dist__q0(krnl_globalSort_L3_0___L4_out_dist__q0),
    .krnl_globalSort_L3_0___L4_out_id__q0(krnl_globalSort_L3_0___L4_out_id__q0),
    .krnl_globalSort_L3_0__ap_start(krnl_globalSort_L3_0__ap_start),
    .krnl_globalSort_L3_0__ap_ready(krnl_globalSort_L3_0__ap_ready),
    .krnl_globalSort_L3_0__ap_done(krnl_globalSort_L3_0__ap_done),
    .krnl_globalSort_L3_0__ap_idle(krnl_globalSort_L3_0__ap_idle),
    .krnl_partialKnn_wrapper_0_0___in_0__q0(krnl_partialKnn_wrapper_0_0___in_0__q0),
    .krnl_partialKnn_wrapper_0_0__ap_start(krnl_partialKnn_wrapper_0_0__ap_start),
    .krnl_partialKnn_wrapper_0_0__ap_ready(krnl_partialKnn_wrapper_0_0__ap_ready),
    .krnl_partialKnn_wrapper_0_0__ap_done(krnl_partialKnn_wrapper_0_0__ap_done),
    .krnl_partialKnn_wrapper_0_0__ap_idle(krnl_partialKnn_wrapper_0_0__ap_idle),
    .krnl_partialKnn_wrapper_1_0___in_1__q0(krnl_partialKnn_wrapper_1_0___in_1__q0),
    .krnl_partialKnn_wrapper_1_0__ap_start(krnl_partialKnn_wrapper_1_0__ap_start),
    .krnl_partialKnn_wrapper_1_0__ap_ready(krnl_partialKnn_wrapper_1_0__ap_ready),
    .krnl_partialKnn_wrapper_1_0__ap_done(krnl_partialKnn_wrapper_1_0__ap_done),
    .krnl_partialKnn_wrapper_1_0__ap_idle(krnl_partialKnn_wrapper_1_0__ap_idle),
    .krnl_partialKnn_wrapper_10_0___in_10__q0(krnl_partialKnn_wrapper_10_0___in_10__q0),
    .krnl_partialKnn_wrapper_10_0__ap_start(krnl_partialKnn_wrapper_10_0__ap_start),
    .krnl_partialKnn_wrapper_10_0__ap_ready(krnl_partialKnn_wrapper_10_0__ap_ready),
    .krnl_partialKnn_wrapper_10_0__ap_done(krnl_partialKnn_wrapper_10_0__ap_done),
    .krnl_partialKnn_wrapper_10_0__ap_idle(krnl_partialKnn_wrapper_10_0__ap_idle),
    .krnl_partialKnn_wrapper_11_0___in_11__q0(krnl_partialKnn_wrapper_11_0___in_11__q0),
    .krnl_partialKnn_wrapper_11_0__ap_start(krnl_partialKnn_wrapper_11_0__ap_start),
    .krnl_partialKnn_wrapper_11_0__ap_ready(krnl_partialKnn_wrapper_11_0__ap_ready),
    .krnl_partialKnn_wrapper_11_0__ap_done(krnl_partialKnn_wrapper_11_0__ap_done),
    .krnl_partialKnn_wrapper_11_0__ap_idle(krnl_partialKnn_wrapper_11_0__ap_idle),
    .krnl_partialKnn_wrapper_12_0___in_12__q0(krnl_partialKnn_wrapper_12_0___in_12__q0),
    .krnl_partialKnn_wrapper_12_0__ap_start(krnl_partialKnn_wrapper_12_0__ap_start),
    .krnl_partialKnn_wrapper_12_0__ap_ready(krnl_partialKnn_wrapper_12_0__ap_ready),
    .krnl_partialKnn_wrapper_12_0__ap_done(krnl_partialKnn_wrapper_12_0__ap_done),
    .krnl_partialKnn_wrapper_12_0__ap_idle(krnl_partialKnn_wrapper_12_0__ap_idle),
    .krnl_partialKnn_wrapper_13_0___in_13__q0(krnl_partialKnn_wrapper_13_0___in_13__q0),
    .krnl_partialKnn_wrapper_13_0__ap_start(krnl_partialKnn_wrapper_13_0__ap_start),
    .krnl_partialKnn_wrapper_13_0__ap_ready(krnl_partialKnn_wrapper_13_0__ap_ready),
    .krnl_partialKnn_wrapper_13_0__ap_done(krnl_partialKnn_wrapper_13_0__ap_done),
    .krnl_partialKnn_wrapper_13_0__ap_idle(krnl_partialKnn_wrapper_13_0__ap_idle),
    .krnl_partialKnn_wrapper_14_0___in_14__q0(krnl_partialKnn_wrapper_14_0___in_14__q0),
    .krnl_partialKnn_wrapper_14_0__ap_start(krnl_partialKnn_wrapper_14_0__ap_start),
    .krnl_partialKnn_wrapper_14_0__ap_ready(krnl_partialKnn_wrapper_14_0__ap_ready),
    .krnl_partialKnn_wrapper_14_0__ap_done(krnl_partialKnn_wrapper_14_0__ap_done),
    .krnl_partialKnn_wrapper_14_0__ap_idle(krnl_partialKnn_wrapper_14_0__ap_idle),
    .krnl_partialKnn_wrapper_15_0___in_15__q0(krnl_partialKnn_wrapper_15_0___in_15__q0),
    .krnl_partialKnn_wrapper_15_0__ap_start(krnl_partialKnn_wrapper_15_0__ap_start),
    .krnl_partialKnn_wrapper_15_0__ap_ready(krnl_partialKnn_wrapper_15_0__ap_ready),
    .krnl_partialKnn_wrapper_15_0__ap_done(krnl_partialKnn_wrapper_15_0__ap_done),
    .krnl_partialKnn_wrapper_15_0__ap_idle(krnl_partialKnn_wrapper_15_0__ap_idle),
    .krnl_partialKnn_wrapper_16_0___in_16__q0(krnl_partialKnn_wrapper_16_0___in_16__q0),
    .krnl_partialKnn_wrapper_16_0__ap_start(krnl_partialKnn_wrapper_16_0__ap_start),
    .krnl_partialKnn_wrapper_16_0__ap_ready(krnl_partialKnn_wrapper_16_0__ap_ready),
    .krnl_partialKnn_wrapper_16_0__ap_done(krnl_partialKnn_wrapper_16_0__ap_done),
    .krnl_partialKnn_wrapper_16_0__ap_idle(krnl_partialKnn_wrapper_16_0__ap_idle),
    .krnl_partialKnn_wrapper_17_0___in_17__q0(krnl_partialKnn_wrapper_17_0___in_17__q0),
    .krnl_partialKnn_wrapper_17_0__ap_start(krnl_partialKnn_wrapper_17_0__ap_start),
    .krnl_partialKnn_wrapper_17_0__ap_ready(krnl_partialKnn_wrapper_17_0__ap_ready),
    .krnl_partialKnn_wrapper_17_0__ap_done(krnl_partialKnn_wrapper_17_0__ap_done),
    .krnl_partialKnn_wrapper_17_0__ap_idle(krnl_partialKnn_wrapper_17_0__ap_idle),
    .krnl_partialKnn_wrapper_18_0___in_18__q0(krnl_partialKnn_wrapper_18_0___in_18__q0),
    .krnl_partialKnn_wrapper_18_0__ap_start(krnl_partialKnn_wrapper_18_0__ap_start),
    .krnl_partialKnn_wrapper_18_0__ap_ready(krnl_partialKnn_wrapper_18_0__ap_ready),
    .krnl_partialKnn_wrapper_18_0__ap_done(krnl_partialKnn_wrapper_18_0__ap_done),
    .krnl_partialKnn_wrapper_18_0__ap_idle(krnl_partialKnn_wrapper_18_0__ap_idle),
    .krnl_partialKnn_wrapper_19_0___in_19__q0(krnl_partialKnn_wrapper_19_0___in_19__q0),
    .krnl_partialKnn_wrapper_19_0__ap_start(krnl_partialKnn_wrapper_19_0__ap_start),
    .krnl_partialKnn_wrapper_19_0__ap_ready(krnl_partialKnn_wrapper_19_0__ap_ready),
    .krnl_partialKnn_wrapper_19_0__ap_done(krnl_partialKnn_wrapper_19_0__ap_done),
    .krnl_partialKnn_wrapper_19_0__ap_idle(krnl_partialKnn_wrapper_19_0__ap_idle),
    .krnl_partialKnn_wrapper_2_0___in_2__q0(krnl_partialKnn_wrapper_2_0___in_2__q0),
    .krnl_partialKnn_wrapper_2_0__ap_start(krnl_partialKnn_wrapper_2_0__ap_start),
    .krnl_partialKnn_wrapper_2_0__ap_ready(krnl_partialKnn_wrapper_2_0__ap_ready),
    .krnl_partialKnn_wrapper_2_0__ap_done(krnl_partialKnn_wrapper_2_0__ap_done),
    .krnl_partialKnn_wrapper_2_0__ap_idle(krnl_partialKnn_wrapper_2_0__ap_idle),
    .krnl_partialKnn_wrapper_20_0___in_20__q0(krnl_partialKnn_wrapper_20_0___in_20__q0),
    .krnl_partialKnn_wrapper_20_0__ap_start(krnl_partialKnn_wrapper_20_0__ap_start),
    .krnl_partialKnn_wrapper_20_0__ap_ready(krnl_partialKnn_wrapper_20_0__ap_ready),
    .krnl_partialKnn_wrapper_20_0__ap_done(krnl_partialKnn_wrapper_20_0__ap_done),
    .krnl_partialKnn_wrapper_20_0__ap_idle(krnl_partialKnn_wrapper_20_0__ap_idle),
    .krnl_partialKnn_wrapper_21_0___in_21__q0(krnl_partialKnn_wrapper_21_0___in_21__q0),
    .krnl_partialKnn_wrapper_21_0__ap_start(krnl_partialKnn_wrapper_21_0__ap_start),
    .krnl_partialKnn_wrapper_21_0__ap_ready(krnl_partialKnn_wrapper_21_0__ap_ready),
    .krnl_partialKnn_wrapper_21_0__ap_done(krnl_partialKnn_wrapper_21_0__ap_done),
    .krnl_partialKnn_wrapper_21_0__ap_idle(krnl_partialKnn_wrapper_21_0__ap_idle),
    .krnl_partialKnn_wrapper_22_0___in_22__q0(krnl_partialKnn_wrapper_22_0___in_22__q0),
    .krnl_partialKnn_wrapper_22_0__ap_start(krnl_partialKnn_wrapper_22_0__ap_start),
    .krnl_partialKnn_wrapper_22_0__ap_ready(krnl_partialKnn_wrapper_22_0__ap_ready),
    .krnl_partialKnn_wrapper_22_0__ap_done(krnl_partialKnn_wrapper_22_0__ap_done),
    .krnl_partialKnn_wrapper_22_0__ap_idle(krnl_partialKnn_wrapper_22_0__ap_idle),
    .krnl_partialKnn_wrapper_23_0___in_23__q0(krnl_partialKnn_wrapper_23_0___in_23__q0),
    .krnl_partialKnn_wrapper_23_0__ap_start(krnl_partialKnn_wrapper_23_0__ap_start),
    .krnl_partialKnn_wrapper_23_0__ap_ready(krnl_partialKnn_wrapper_23_0__ap_ready),
    .krnl_partialKnn_wrapper_23_0__ap_done(krnl_partialKnn_wrapper_23_0__ap_done),
    .krnl_partialKnn_wrapper_23_0__ap_idle(krnl_partialKnn_wrapper_23_0__ap_idle),
    .krnl_partialKnn_wrapper_24_0___in_24__q0(krnl_partialKnn_wrapper_24_0___in_24__q0),
    .krnl_partialKnn_wrapper_24_0__ap_start(krnl_partialKnn_wrapper_24_0__ap_start),
    .krnl_partialKnn_wrapper_24_0__ap_ready(krnl_partialKnn_wrapper_24_0__ap_ready),
    .krnl_partialKnn_wrapper_24_0__ap_done(krnl_partialKnn_wrapper_24_0__ap_done),
    .krnl_partialKnn_wrapper_24_0__ap_idle(krnl_partialKnn_wrapper_24_0__ap_idle),
    .krnl_partialKnn_wrapper_25_0___in_25__q0(krnl_partialKnn_wrapper_25_0___in_25__q0),
    .krnl_partialKnn_wrapper_25_0__ap_start(krnl_partialKnn_wrapper_25_0__ap_start),
    .krnl_partialKnn_wrapper_25_0__ap_ready(krnl_partialKnn_wrapper_25_0__ap_ready),
    .krnl_partialKnn_wrapper_25_0__ap_done(krnl_partialKnn_wrapper_25_0__ap_done),
    .krnl_partialKnn_wrapper_25_0__ap_idle(krnl_partialKnn_wrapper_25_0__ap_idle),
    .krnl_partialKnn_wrapper_26_0___in_26__q0(krnl_partialKnn_wrapper_26_0___in_26__q0),
    .krnl_partialKnn_wrapper_26_0__ap_start(krnl_partialKnn_wrapper_26_0__ap_start),
    .krnl_partialKnn_wrapper_26_0__ap_ready(krnl_partialKnn_wrapper_26_0__ap_ready),
    .krnl_partialKnn_wrapper_26_0__ap_done(krnl_partialKnn_wrapper_26_0__ap_done),
    .krnl_partialKnn_wrapper_26_0__ap_idle(krnl_partialKnn_wrapper_26_0__ap_idle),
    .krnl_partialKnn_wrapper_27_0___in_27__q0(krnl_partialKnn_wrapper_27_0___in_27__q0),
    .krnl_partialKnn_wrapper_27_0__ap_start(krnl_partialKnn_wrapper_27_0__ap_start),
    .krnl_partialKnn_wrapper_27_0__ap_ready(krnl_partialKnn_wrapper_27_0__ap_ready),
    .krnl_partialKnn_wrapper_27_0__ap_done(krnl_partialKnn_wrapper_27_0__ap_done),
    .krnl_partialKnn_wrapper_27_0__ap_idle(krnl_partialKnn_wrapper_27_0__ap_idle),
    .krnl_partialKnn_wrapper_28_0___in_28__q0(krnl_partialKnn_wrapper_28_0___in_28__q0),
    .krnl_partialKnn_wrapper_28_0__ap_start(krnl_partialKnn_wrapper_28_0__ap_start),
    .krnl_partialKnn_wrapper_28_0__ap_ready(krnl_partialKnn_wrapper_28_0__ap_ready),
    .krnl_partialKnn_wrapper_28_0__ap_done(krnl_partialKnn_wrapper_28_0__ap_done),
    .krnl_partialKnn_wrapper_28_0__ap_idle(krnl_partialKnn_wrapper_28_0__ap_idle),
    .krnl_partialKnn_wrapper_29_0___in_29__q0(krnl_partialKnn_wrapper_29_0___in_29__q0),
    .krnl_partialKnn_wrapper_29_0__ap_start(krnl_partialKnn_wrapper_29_0__ap_start),
    .krnl_partialKnn_wrapper_29_0__ap_ready(krnl_partialKnn_wrapper_29_0__ap_ready),
    .krnl_partialKnn_wrapper_29_0__ap_done(krnl_partialKnn_wrapper_29_0__ap_done),
    .krnl_partialKnn_wrapper_29_0__ap_idle(krnl_partialKnn_wrapper_29_0__ap_idle),
    .krnl_partialKnn_wrapper_3_0___in_3__q0(krnl_partialKnn_wrapper_3_0___in_3__q0),
    .krnl_partialKnn_wrapper_3_0__ap_start(krnl_partialKnn_wrapper_3_0__ap_start),
    .krnl_partialKnn_wrapper_3_0__ap_ready(krnl_partialKnn_wrapper_3_0__ap_ready),
    .krnl_partialKnn_wrapper_3_0__ap_done(krnl_partialKnn_wrapper_3_0__ap_done),
    .krnl_partialKnn_wrapper_3_0__ap_idle(krnl_partialKnn_wrapper_3_0__ap_idle),
    .krnl_partialKnn_wrapper_30_0___in_30__q0(krnl_partialKnn_wrapper_30_0___in_30__q0),
    .krnl_partialKnn_wrapper_30_0__ap_start(krnl_partialKnn_wrapper_30_0__ap_start),
    .krnl_partialKnn_wrapper_30_0__ap_ready(krnl_partialKnn_wrapper_30_0__ap_ready),
    .krnl_partialKnn_wrapper_30_0__ap_done(krnl_partialKnn_wrapper_30_0__ap_done),
    .krnl_partialKnn_wrapper_30_0__ap_idle(krnl_partialKnn_wrapper_30_0__ap_idle),
    .krnl_partialKnn_wrapper_31_0___in_31__q0(krnl_partialKnn_wrapper_31_0___in_31__q0),
    .krnl_partialKnn_wrapper_31_0__ap_start(krnl_partialKnn_wrapper_31_0__ap_start),
    .krnl_partialKnn_wrapper_31_0__ap_ready(krnl_partialKnn_wrapper_31_0__ap_ready),
    .krnl_partialKnn_wrapper_31_0__ap_done(krnl_partialKnn_wrapper_31_0__ap_done),
    .krnl_partialKnn_wrapper_31_0__ap_idle(krnl_partialKnn_wrapper_31_0__ap_idle),
    .krnl_partialKnn_wrapper_32_0___in_32__q0(krnl_partialKnn_wrapper_32_0___in_32__q0),
    .krnl_partialKnn_wrapper_32_0__ap_start(krnl_partialKnn_wrapper_32_0__ap_start),
    .krnl_partialKnn_wrapper_32_0__ap_ready(krnl_partialKnn_wrapper_32_0__ap_ready),
    .krnl_partialKnn_wrapper_32_0__ap_done(krnl_partialKnn_wrapper_32_0__ap_done),
    .krnl_partialKnn_wrapper_32_0__ap_idle(krnl_partialKnn_wrapper_32_0__ap_idle),
    .krnl_partialKnn_wrapper_33_0___in_33__q0(krnl_partialKnn_wrapper_33_0___in_33__q0),
    .krnl_partialKnn_wrapper_33_0__ap_start(krnl_partialKnn_wrapper_33_0__ap_start),
    .krnl_partialKnn_wrapper_33_0__ap_ready(krnl_partialKnn_wrapper_33_0__ap_ready),
    .krnl_partialKnn_wrapper_33_0__ap_done(krnl_partialKnn_wrapper_33_0__ap_done),
    .krnl_partialKnn_wrapper_33_0__ap_idle(krnl_partialKnn_wrapper_33_0__ap_idle),
    .krnl_partialKnn_wrapper_34_0___in_34__q0(krnl_partialKnn_wrapper_34_0___in_34__q0),
    .krnl_partialKnn_wrapper_34_0__ap_start(krnl_partialKnn_wrapper_34_0__ap_start),
    .krnl_partialKnn_wrapper_34_0__ap_ready(krnl_partialKnn_wrapper_34_0__ap_ready),
    .krnl_partialKnn_wrapper_34_0__ap_done(krnl_partialKnn_wrapper_34_0__ap_done),
    .krnl_partialKnn_wrapper_34_0__ap_idle(krnl_partialKnn_wrapper_34_0__ap_idle),
    .krnl_partialKnn_wrapper_35_0___in_35__q0(krnl_partialKnn_wrapper_35_0___in_35__q0),
    .krnl_partialKnn_wrapper_35_0__ap_start(krnl_partialKnn_wrapper_35_0__ap_start),
    .krnl_partialKnn_wrapper_35_0__ap_ready(krnl_partialKnn_wrapper_35_0__ap_ready),
    .krnl_partialKnn_wrapper_35_0__ap_done(krnl_partialKnn_wrapper_35_0__ap_done),
    .krnl_partialKnn_wrapper_35_0__ap_idle(krnl_partialKnn_wrapper_35_0__ap_idle),
    .krnl_partialKnn_wrapper_36_0___in_36__q0(krnl_partialKnn_wrapper_36_0___in_36__q0),
    .krnl_partialKnn_wrapper_36_0__ap_start(krnl_partialKnn_wrapper_36_0__ap_start),
    .krnl_partialKnn_wrapper_36_0__ap_ready(krnl_partialKnn_wrapper_36_0__ap_ready),
    .krnl_partialKnn_wrapper_36_0__ap_done(krnl_partialKnn_wrapper_36_0__ap_done),
    .krnl_partialKnn_wrapper_36_0__ap_idle(krnl_partialKnn_wrapper_36_0__ap_idle),
    .krnl_partialKnn_wrapper_37_0___in_37__q0(krnl_partialKnn_wrapper_37_0___in_37__q0),
    .krnl_partialKnn_wrapper_37_0__ap_start(krnl_partialKnn_wrapper_37_0__ap_start),
    .krnl_partialKnn_wrapper_37_0__ap_ready(krnl_partialKnn_wrapper_37_0__ap_ready),
    .krnl_partialKnn_wrapper_37_0__ap_done(krnl_partialKnn_wrapper_37_0__ap_done),
    .krnl_partialKnn_wrapper_37_0__ap_idle(krnl_partialKnn_wrapper_37_0__ap_idle),
    .krnl_partialKnn_wrapper_38_0___in_38__q0(krnl_partialKnn_wrapper_38_0___in_38__q0),
    .krnl_partialKnn_wrapper_38_0__ap_start(krnl_partialKnn_wrapper_38_0__ap_start),
    .krnl_partialKnn_wrapper_38_0__ap_ready(krnl_partialKnn_wrapper_38_0__ap_ready),
    .krnl_partialKnn_wrapper_38_0__ap_done(krnl_partialKnn_wrapper_38_0__ap_done),
    .krnl_partialKnn_wrapper_38_0__ap_idle(krnl_partialKnn_wrapper_38_0__ap_idle),
    .krnl_partialKnn_wrapper_39_0___in_39__q0(krnl_partialKnn_wrapper_39_0___in_39__q0),
    .krnl_partialKnn_wrapper_39_0__ap_start(krnl_partialKnn_wrapper_39_0__ap_start),
    .krnl_partialKnn_wrapper_39_0__ap_ready(krnl_partialKnn_wrapper_39_0__ap_ready),
    .krnl_partialKnn_wrapper_39_0__ap_done(krnl_partialKnn_wrapper_39_0__ap_done),
    .krnl_partialKnn_wrapper_39_0__ap_idle(krnl_partialKnn_wrapper_39_0__ap_idle),
    .krnl_partialKnn_wrapper_4_0___in_4__q0(krnl_partialKnn_wrapper_4_0___in_4__q0),
    .krnl_partialKnn_wrapper_4_0__ap_start(krnl_partialKnn_wrapper_4_0__ap_start),
    .krnl_partialKnn_wrapper_4_0__ap_ready(krnl_partialKnn_wrapper_4_0__ap_ready),
    .krnl_partialKnn_wrapper_4_0__ap_done(krnl_partialKnn_wrapper_4_0__ap_done),
    .krnl_partialKnn_wrapper_4_0__ap_idle(krnl_partialKnn_wrapper_4_0__ap_idle),
    .krnl_partialKnn_wrapper_40_0___in_40__q0(krnl_partialKnn_wrapper_40_0___in_40__q0),
    .krnl_partialKnn_wrapper_40_0__ap_start(krnl_partialKnn_wrapper_40_0__ap_start),
    .krnl_partialKnn_wrapper_40_0__ap_ready(krnl_partialKnn_wrapper_40_0__ap_ready),
    .krnl_partialKnn_wrapper_40_0__ap_done(krnl_partialKnn_wrapper_40_0__ap_done),
    .krnl_partialKnn_wrapper_40_0__ap_idle(krnl_partialKnn_wrapper_40_0__ap_idle),
    .krnl_partialKnn_wrapper_41_0___in_41__q0(krnl_partialKnn_wrapper_41_0___in_41__q0),
    .krnl_partialKnn_wrapper_41_0__ap_start(krnl_partialKnn_wrapper_41_0__ap_start),
    .krnl_partialKnn_wrapper_41_0__ap_ready(krnl_partialKnn_wrapper_41_0__ap_ready),
    .krnl_partialKnn_wrapper_41_0__ap_done(krnl_partialKnn_wrapper_41_0__ap_done),
    .krnl_partialKnn_wrapper_41_0__ap_idle(krnl_partialKnn_wrapper_41_0__ap_idle),
    .krnl_partialKnn_wrapper_42_0___in_42__q0(krnl_partialKnn_wrapper_42_0___in_42__q0),
    .krnl_partialKnn_wrapper_42_0__ap_start(krnl_partialKnn_wrapper_42_0__ap_start),
    .krnl_partialKnn_wrapper_42_0__ap_ready(krnl_partialKnn_wrapper_42_0__ap_ready),
    .krnl_partialKnn_wrapper_42_0__ap_done(krnl_partialKnn_wrapper_42_0__ap_done),
    .krnl_partialKnn_wrapper_42_0__ap_idle(krnl_partialKnn_wrapper_42_0__ap_idle),
    .krnl_partialKnn_wrapper_43_0___in_43__q0(krnl_partialKnn_wrapper_43_0___in_43__q0),
    .krnl_partialKnn_wrapper_43_0__ap_start(krnl_partialKnn_wrapper_43_0__ap_start),
    .krnl_partialKnn_wrapper_43_0__ap_ready(krnl_partialKnn_wrapper_43_0__ap_ready),
    .krnl_partialKnn_wrapper_43_0__ap_done(krnl_partialKnn_wrapper_43_0__ap_done),
    .krnl_partialKnn_wrapper_43_0__ap_idle(krnl_partialKnn_wrapper_43_0__ap_idle),
    .krnl_partialKnn_wrapper_44_0___in_44__q0(krnl_partialKnn_wrapper_44_0___in_44__q0),
    .krnl_partialKnn_wrapper_44_0__ap_start(krnl_partialKnn_wrapper_44_0__ap_start),
    .krnl_partialKnn_wrapper_44_0__ap_ready(krnl_partialKnn_wrapper_44_0__ap_ready),
    .krnl_partialKnn_wrapper_44_0__ap_done(krnl_partialKnn_wrapper_44_0__ap_done),
    .krnl_partialKnn_wrapper_44_0__ap_idle(krnl_partialKnn_wrapper_44_0__ap_idle),
    .krnl_partialKnn_wrapper_45_0___in_45__q0(krnl_partialKnn_wrapper_45_0___in_45__q0),
    .krnl_partialKnn_wrapper_45_0__ap_start(krnl_partialKnn_wrapper_45_0__ap_start),
    .krnl_partialKnn_wrapper_45_0__ap_ready(krnl_partialKnn_wrapper_45_0__ap_ready),
    .krnl_partialKnn_wrapper_45_0__ap_done(krnl_partialKnn_wrapper_45_0__ap_done),
    .krnl_partialKnn_wrapper_45_0__ap_idle(krnl_partialKnn_wrapper_45_0__ap_idle),
    .krnl_partialKnn_wrapper_46_0___in_46__q0(krnl_partialKnn_wrapper_46_0___in_46__q0),
    .krnl_partialKnn_wrapper_46_0__ap_start(krnl_partialKnn_wrapper_46_0__ap_start),
    .krnl_partialKnn_wrapper_46_0__ap_ready(krnl_partialKnn_wrapper_46_0__ap_ready),
    .krnl_partialKnn_wrapper_46_0__ap_done(krnl_partialKnn_wrapper_46_0__ap_done),
    .krnl_partialKnn_wrapper_46_0__ap_idle(krnl_partialKnn_wrapper_46_0__ap_idle),
    .krnl_partialKnn_wrapper_47_0___in_47__q0(krnl_partialKnn_wrapper_47_0___in_47__q0),
    .krnl_partialKnn_wrapper_47_0__ap_start(krnl_partialKnn_wrapper_47_0__ap_start),
    .krnl_partialKnn_wrapper_47_0__ap_ready(krnl_partialKnn_wrapper_47_0__ap_ready),
    .krnl_partialKnn_wrapper_47_0__ap_done(krnl_partialKnn_wrapper_47_0__ap_done),
    .krnl_partialKnn_wrapper_47_0__ap_idle(krnl_partialKnn_wrapper_47_0__ap_idle),
    .krnl_partialKnn_wrapper_48_0___in_48__q0(krnl_partialKnn_wrapper_48_0___in_48__q0),
    .krnl_partialKnn_wrapper_48_0__ap_start(krnl_partialKnn_wrapper_48_0__ap_start),
    .krnl_partialKnn_wrapper_48_0__ap_ready(krnl_partialKnn_wrapper_48_0__ap_ready),
    .krnl_partialKnn_wrapper_48_0__ap_done(krnl_partialKnn_wrapper_48_0__ap_done),
    .krnl_partialKnn_wrapper_48_0__ap_idle(krnl_partialKnn_wrapper_48_0__ap_idle),
    .krnl_partialKnn_wrapper_49_0___in_49__q0(krnl_partialKnn_wrapper_49_0___in_49__q0),
    .krnl_partialKnn_wrapper_49_0__ap_start(krnl_partialKnn_wrapper_49_0__ap_start),
    .krnl_partialKnn_wrapper_49_0__ap_ready(krnl_partialKnn_wrapper_49_0__ap_ready),
    .krnl_partialKnn_wrapper_49_0__ap_done(krnl_partialKnn_wrapper_49_0__ap_done),
    .krnl_partialKnn_wrapper_49_0__ap_idle(krnl_partialKnn_wrapper_49_0__ap_idle),
    .krnl_partialKnn_wrapper_5_0___in_5__q0(krnl_partialKnn_wrapper_5_0___in_5__q0),
    .krnl_partialKnn_wrapper_5_0__ap_start(krnl_partialKnn_wrapper_5_0__ap_start),
    .krnl_partialKnn_wrapper_5_0__ap_ready(krnl_partialKnn_wrapper_5_0__ap_ready),
    .krnl_partialKnn_wrapper_5_0__ap_done(krnl_partialKnn_wrapper_5_0__ap_done),
    .krnl_partialKnn_wrapper_5_0__ap_idle(krnl_partialKnn_wrapper_5_0__ap_idle),
    .krnl_partialKnn_wrapper_50_0___in_50__q0(krnl_partialKnn_wrapper_50_0___in_50__q0),
    .krnl_partialKnn_wrapper_50_0__ap_start(krnl_partialKnn_wrapper_50_0__ap_start),
    .krnl_partialKnn_wrapper_50_0__ap_ready(krnl_partialKnn_wrapper_50_0__ap_ready),
    .krnl_partialKnn_wrapper_50_0__ap_done(krnl_partialKnn_wrapper_50_0__ap_done),
    .krnl_partialKnn_wrapper_50_0__ap_idle(krnl_partialKnn_wrapper_50_0__ap_idle),
    .krnl_partialKnn_wrapper_51_0___in_51__q0(krnl_partialKnn_wrapper_51_0___in_51__q0),
    .krnl_partialKnn_wrapper_51_0__ap_start(krnl_partialKnn_wrapper_51_0__ap_start),
    .krnl_partialKnn_wrapper_51_0__ap_ready(krnl_partialKnn_wrapper_51_0__ap_ready),
    .krnl_partialKnn_wrapper_51_0__ap_done(krnl_partialKnn_wrapper_51_0__ap_done),
    .krnl_partialKnn_wrapper_51_0__ap_idle(krnl_partialKnn_wrapper_51_0__ap_idle),
    .krnl_partialKnn_wrapper_52_0___in_52__q0(krnl_partialKnn_wrapper_52_0___in_52__q0),
    .krnl_partialKnn_wrapper_52_0__ap_start(krnl_partialKnn_wrapper_52_0__ap_start),
    .krnl_partialKnn_wrapper_52_0__ap_ready(krnl_partialKnn_wrapper_52_0__ap_ready),
    .krnl_partialKnn_wrapper_52_0__ap_done(krnl_partialKnn_wrapper_52_0__ap_done),
    .krnl_partialKnn_wrapper_52_0__ap_idle(krnl_partialKnn_wrapper_52_0__ap_idle),
    .krnl_partialKnn_wrapper_53_0___in_53__q0(krnl_partialKnn_wrapper_53_0___in_53__q0),
    .krnl_partialKnn_wrapper_53_0__ap_start(krnl_partialKnn_wrapper_53_0__ap_start),
    .krnl_partialKnn_wrapper_53_0__ap_ready(krnl_partialKnn_wrapper_53_0__ap_ready),
    .krnl_partialKnn_wrapper_53_0__ap_done(krnl_partialKnn_wrapper_53_0__ap_done),
    .krnl_partialKnn_wrapper_53_0__ap_idle(krnl_partialKnn_wrapper_53_0__ap_idle),
    .krnl_partialKnn_wrapper_6_0___in_6__q0(krnl_partialKnn_wrapper_6_0___in_6__q0),
    .krnl_partialKnn_wrapper_6_0__ap_start(krnl_partialKnn_wrapper_6_0__ap_start),
    .krnl_partialKnn_wrapper_6_0__ap_ready(krnl_partialKnn_wrapper_6_0__ap_ready),
    .krnl_partialKnn_wrapper_6_0__ap_done(krnl_partialKnn_wrapper_6_0__ap_done),
    .krnl_partialKnn_wrapper_6_0__ap_idle(krnl_partialKnn_wrapper_6_0__ap_idle),
    .krnl_partialKnn_wrapper_7_0___in_7__q0(krnl_partialKnn_wrapper_7_0___in_7__q0),
    .krnl_partialKnn_wrapper_7_0__ap_start(krnl_partialKnn_wrapper_7_0__ap_start),
    .krnl_partialKnn_wrapper_7_0__ap_ready(krnl_partialKnn_wrapper_7_0__ap_ready),
    .krnl_partialKnn_wrapper_7_0__ap_done(krnl_partialKnn_wrapper_7_0__ap_done),
    .krnl_partialKnn_wrapper_7_0__ap_idle(krnl_partialKnn_wrapper_7_0__ap_idle),
    .krnl_partialKnn_wrapper_8_0___in_8__q0(krnl_partialKnn_wrapper_8_0___in_8__q0),
    .krnl_partialKnn_wrapper_8_0__ap_start(krnl_partialKnn_wrapper_8_0__ap_start),
    .krnl_partialKnn_wrapper_8_0__ap_ready(krnl_partialKnn_wrapper_8_0__ap_ready),
    .krnl_partialKnn_wrapper_8_0__ap_done(krnl_partialKnn_wrapper_8_0__ap_done),
    .krnl_partialKnn_wrapper_8_0__ap_idle(krnl_partialKnn_wrapper_8_0__ap_idle),
    .krnl_partialKnn_wrapper_9_0___in_9__q0(krnl_partialKnn_wrapper_9_0___in_9__q0),
    .krnl_partialKnn_wrapper_9_0__ap_start(krnl_partialKnn_wrapper_9_0__ap_start),
    .krnl_partialKnn_wrapper_9_0__ap_ready(krnl_partialKnn_wrapper_9_0__ap_ready),
    .krnl_partialKnn_wrapper_9_0__ap_done(krnl_partialKnn_wrapper_9_0__ap_done),
    .krnl_partialKnn_wrapper_9_0__ap_idle(krnl_partialKnn_wrapper_9_0__ap_idle)
  );

  assign ap_rst_n_inv = (~ap_rst_n);

endmodule

